----------------------------------------------------------------------
-- Created by Actel SmartDesign Thu Apr 23 15:24:11 2009
-- Parameters for COREUART
----------------------------------------------------------------------


package coreparameters is
    constant FAMILY : integer := 20;
    constant HDL_license : string( 1 to 1 ) := "O";
    constant RX_FIFO : integer := 0;
    constant TX_FIFO : integer := 0;
    constant testbench : string( 1 to 5 ) := "Verif";
end coreparameters;
