-- Rev:			2.2 24Jan05 TFB - Production


library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity XYXX0008 is

   port( XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0 : in std_logic;  
         XXXXXXXXXXXXXXXXXJXXXXX : out std_logic;  XLX, XXXXXXXX : in std_logic
         ;  JXXXXX, XXXXXX : out std_logic;  
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX : in std_logic;  XXXXXXXX0 : 
         out std_logic;  MXMXXXXXXXX : in std_logic;  MXMXXXX : in 
         std_logic_vector (15 downto 0);  XXXXXXX : in std_logic_vector (19 
         downto 0);  XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXPX, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, XXXXXXXX1, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXP, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH : in std_logic;  MXMXXXX0 : 
         in std_logic_vector (3 downto 0);  MXMXXXXXXXX0, XXXXXXXX2, 
         MXMXXXXXXXX1, MXMXXXXXXXX2, XXXXXXXX3, XXXXXXXX4, XXXXXXXX5 : in 
         std_logic;  XXXXXXXXP : out std_logic;  
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX1, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX2, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX3, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX4, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX5, 
         XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX6, XXXXXX0 : in std_logic; 
         XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, 
         XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, 
         XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1, 
         XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2, 
         XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3, 
         XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4, 
         XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5, 
         XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6 : out std_logic;  XXXXXXXX6
         , XXXXXXXX7 : in std_logic;  XXXXXPXWX, XXXXXPXXX, XXXXXXXX8 : out 
         std_logic;  XXXXXXX0, XXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXX, MXMPXXXXX : 
         in std_logic);

end XYXX0008;

architecture SYN_USE_DEFA_ARCH_NAME of XYXX0008 is

signal XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXLXXXXXX, XXXXXXXXXXXXXXXXXJXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, XXXXXXXXXXXXXXXXXXXXXX, 
   XXXXXXXXXXXXXXXXXJXXXXX1, XXXXXXXXXXXXXXXXXXXXXX0, XXXXXXXXXXXXXXXXXJXXXXX2,
   XXXXXXXXXXXXXXXXXXXXXX1, XXXXXXXXXXXXXXXXXJXXXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX11, XXXXXXXXXXXXXXXXXJXXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, XXXXXXXXXXXXXXXXXJXXXXX5, 
   XXXXXXXXXXXXXXXXXXXXXX2, XXXXXXXXXXXXXXXXXJXXXXX6, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3, XXXXXXXXXXXXXXXXXXXXXX3, 
   XXXXXXXXXXXXXXXXXJXXXXX7, XXXXXXXXXXXXXXXXXXXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX29, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX5, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX30, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX6, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX31, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX7, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX32, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX8, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX33, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX9, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX34, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX10, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX35, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX11, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX36, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX12, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX37, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX13, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX38, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX14, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX39, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX15, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX40, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX16, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX41, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX17, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX42, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX18, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX43, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX19, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX44, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX20, XXXXXXXXXXXXXXXXXJXXXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX21, XXXXXXXXXXXXXXXXXJXXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX22, XXXXXXXXXXXXXXXXXJXXXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX23, XXXXXXXXXXXXXXXXXJXXXXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX24, XXXXXXXXXXXXXXXXXJXXXXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX25, XXXXXXXXXXXXXXXXXJXXXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX26, XXXXXXXXXXXXXXXXXJXXXXXX5, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX27, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, XXXXXXXXXXXXXXXXXJXXXXXX6, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX28, XXXXXXXXXXXXXXXXXJXXXXXX7, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX29, XXXXXXXXXXXXXXXXXJXXXXXX8, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX30, XXXXXXXXXXXXXXXXXJXXXXXX9, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX31, XXXXXXXXXXXXXXXXXJXXXXXX10, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX32, XXXXXXXXXXXXXXXXXJXXXXXX11, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX33, XXXXXXXXXXXXXXXXXJXXXXXX12, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX10, XXXXXXXXXXXXXXXXXJXXXXX8, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX11, XXXXXXXXXXXXXXXXXJXXXXX9, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX12, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX13, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX14, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX15, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX16, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX17, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX18, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX19, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXXXHXLXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXYXXXXXXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX5, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX6, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX34, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX, XXXXXXXXXXXXXXXXXJXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX0, XXXXXXXXXXXXXXXXXJXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXYXXXXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX20, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX21, XXXXXXXX00, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX7, XXXXXXXXXXXXXXXXXXXXXXXXXYPX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX8, XXXXXXXXXXXXXXXXXXXXXXXXXYPX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX9, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX10, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX22, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXMXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX23, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX24, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX25, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX26, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX4, 
   XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX35, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX29, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX30, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX31, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX12, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXJXXXXXHXLXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX36, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX37, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX38, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX39, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX40, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX41, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX42, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX43, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX44, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX45, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX32, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX33, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX5, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX6, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX7, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX8, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX9, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX10, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX11, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX12, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX13, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX46, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX5, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX6, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX7, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX8, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX9, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX10, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX11, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX12, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX13, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXXXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX0, XXXXXXXXXXXXXXXXXXXXXX5, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX11, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX5, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX6, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX1, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX5, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX6, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX7, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX8, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX9, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX16, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX10, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX7, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX8, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX12, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX9, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX10, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX11, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX12, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX13, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX14, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX15, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX16, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX17, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX18, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX19, XXXXXXXXP0, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX20, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXXXX, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX2, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX21, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX3, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX22, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX4, 
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX23, 
   XXXXXXXXXXXXXXXXXXXXXXXX, XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX15, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX0, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX00, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX1, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX16, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX2, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX20, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX3, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX30, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX4, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX40, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX5, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX50, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX6, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX60, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX7, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX23, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX8, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX24, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX9, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX25, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX10, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX26, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX11, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX27, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX12, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX28, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX0, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX0, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX1, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX2, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX3, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX4, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX5, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX6, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX7, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX8, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX0, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXYPXXXHXL, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXLXY, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXL, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXHXLXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXX0, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXPXXHXLXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXMXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXXHXL, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX13, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXX0, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX14, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXYPXXXHXLXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX15, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX16, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX17, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX18, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX19, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX20, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX21, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX22, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX23, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX24, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX25, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX26, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX1, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX2, 
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX0
   : std_logic;

begin
   XXXXXXXXXXXXXXXXXJXXXXX <= XXXXXXXXXXXXXXXXXJXXXXX7;
   XXXXXXXX0 <= XXXXXXXX00;
   XXXXXXXXP <= XXXXXXXXP0;
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX <= 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX15;
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0 <= 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX00;
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1 <= 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX16;
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2 <= 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX20;
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3 <= 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX30;
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4 <= 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX40;
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5 <= 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX50;
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6 <= 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX60;
   
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXLXXXXXX <= '0';
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX0, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX1, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX2, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX4 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX3, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX11);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX5 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX4, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX6 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX5, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXXXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX7 : DFN1E1P0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX6, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, PRE => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXXXXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX8 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX7, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXXXXXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX4, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX29);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX0 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX5, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX30);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX1 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX6, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX31);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX2 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX7, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX32);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX3 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX8, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX33);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX4 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX9, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX34);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX5 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX10, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX35);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX6 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX11, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX36);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX7 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX12, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX37);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX8 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX13, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX38);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX9 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX14, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX39);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX10 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX15, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX40);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX11 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX16, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX41);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX12 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX17, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX42);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX13 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX18, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX43);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX14 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX19, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX44);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX15 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX20, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX16 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX21, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX17 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX22, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX18 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX23, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX19 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX24, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX20 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX25, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX21 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX26, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX5);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX22 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX27, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX6);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX23 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX28, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX7);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX24 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX29, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX8);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX25 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX30, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX9);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX26 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX31, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX10);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX27 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX32, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX11);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX28 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX33, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXXX12);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX10, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX8);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX0 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX11, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX9);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX1 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX12, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX2 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX13, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX3 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX14, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX4 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX15, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX5 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX16, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX6 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX17, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX5);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX7 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX18, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX6);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX8 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX19, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXJXXXXX7);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXXXXXXX : DFN1P0 port map( D
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXXXXXX, 
                           CLK => XLX, PRE => XXXXXXXX, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXX0)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXX9 : DFN1E0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXXXHXLXX, E 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXYXXXXXXXXX, 
                           CLK => XLX, Q => JXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX6, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPX0, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX5, CLK => 
                           XLX, CLR => XXXXXXXX, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX6, CLK => 
                           XLX, CLR => XXXXXXXX, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX5);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX34, CLK 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX6);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXX : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX, CLK 
                           => XLX, CLR => XXXXXXXX, Q => XXXXXXXXXXXXXXXXXJXXX)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXX0 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX0, CLK 
                           => XLX, CLR => XXXXXXXX, Q => XXXXXXXXXXXXXXXXXJXXX0
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXYXXXXXXXXXXXX : DFN1P0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXLXXXXXX, CLK => 
                           XLX, PRE => XXXXXXXX, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXYXXXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX1 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX0, CLK => XLX
                           , CLR => XXXXXXXX, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX1, CLK => XLX
                           , CLR => XXXXXXXX, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX7 : NOR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX2, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX8 : NOR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX9 : MX2C port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX6, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX20, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX9, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX21);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX1 : MX2 port map( A => 
                           XXXXXXXX00, S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX4, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX7);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX2 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXXXXXYPX, S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX1, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX8);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX3 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXXXXXYPX0, S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX9);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX4 : OR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX7, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX10);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXXXXXXX : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX, B =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX10, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXX : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXX4, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXXXXXX : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX22, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXMXXXXXXXX : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX1, B 
                           => MXMXXXXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXMXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXXXXXX0 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX23, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXXXXXX1 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX24, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXXXXXX2 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX21, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX2, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX23);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX0 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX0 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX1, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX22);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX44, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX1 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX43, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX, Y =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX19);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX1 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX30, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX2 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX31, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX1, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX6);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           MXMXXXX(0), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(0), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX25);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX1 : MX2 port map( A => 
                           MXMXXXX(3), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(3), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX22);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX2 : MX2 port map( A => 
                           MXMXXXX(5), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(5), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX23);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX3 : MX2 port map( A => 
                           MXMXXXX(6), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(6), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX24);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX4 : MX2 port map( A => 
                           MXMXXXX(7), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(7), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX26);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX0 : OR3 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX3, 
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, Y
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX5 : OR2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX, B =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX4, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXXXHXLXXXXXXX : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX11, S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXYXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXXXHXLXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXYXXXXXXXXXXXXXX : NOR2A port map( A 
                           => XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXYXXXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXYXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXX0,
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXXXXXXX : OR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXXXXX0, C => XXXXXXXXXXXXXXXXXXXXXX
                           , Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX1 : NOR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX0, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXPX, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX34);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPX : NOR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX1, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXPX, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX : MX2C port map( A => XXXXXXXX1, 
                           S => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, 
                           B => XXXXXXXXXXXXXXXXXJXXXXX5, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX35);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXX0 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXX2, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX5 : MX2 port map( A => 
                           MXMXXXX(2), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(2), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX29);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX6 : MX2 port map( A => 
                           MXMXXXX(4), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(4), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX30);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX7 : MX2 port map( A => 
                           MXMXXXX(1), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(1), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX31);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXXXXXX3 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX31, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX6 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXX0,
                           S => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, 
                           B => XXXXXXXXXXXXXXXXXJXXXXX6, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX12);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXJXXXXXHXL : AO16 port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXXXXX1, C => XXXXXXXXXXXXXXXXXXXXXX
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXJXXXXXHXLXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXXXXX : OR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX1, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXP, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXXXXX0 : NOR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX0, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXP, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXX : NOR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX1, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXX0 : NOR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX0, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX0 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX29, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX2 : MX2 port map( A => 
                           MXMXXXX0(3), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(19), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX36);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX3 : MX2 port map( A => 
                           MXMXXXX0(2), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX12, B => 
                           XXXXXXX(18), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX37);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX4 : MX2 port map( A => 
                           MXMXXXX0(1), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(17), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX38);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX5 : MX2 port map( A => 
                           MXMXXXX0(0), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(16), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX39);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX6 : MX2 port map( A => 
                           MXMXXXX(15), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(15), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX40);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX7 : MX2 port map( A => 
                           MXMXXXX(14), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(14), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX41);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX8 : MX2 port map( A => 
                           MXMXXXX(13), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(13), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX42);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX9 : MX2 port map( A => 
                           MXMXXXX(12), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(12), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX43);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX10 : MX2 port map( A => 
                           MXMXXXX(11), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(11), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX44);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX11 : MX2 port map( A => 
                           MXMXXXX(10), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(10), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX45);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX8 : MX2 port map( A => 
                           MXMXXXX(9), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(9), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX32);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX9 : MX2 port map( A => 
                           MXMXXXX(8), S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, B => 
                           XXXXXXX(8), Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX33);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX3 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX29, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX1, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX5);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX1 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX30, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX4 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX31, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX2, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX7);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX2 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX32, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX5 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX32, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX3, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX8);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX3 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX33, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX6 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX33, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX4, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX9);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX4 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX34, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX7 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX34, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX5, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX10);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX5 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX35, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX5);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX8 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX13, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX35, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX6, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX11);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX6 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX36, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX6);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX9 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX36, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX7, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX12);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX7 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX37, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX7);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX10 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX37, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX8, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX13);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX8 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX38, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX8);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX11 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX38, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX9, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX14);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX9 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX39, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX9);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX12 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX39, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX10, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX15);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX10 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX40, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX10);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX13 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX40, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX11, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX16);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX11 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX41, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX11);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX14 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX41, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX12, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX17);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX12 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX42, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX12);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX15 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX42, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX13, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX18);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXXXX13 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX43, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX13);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXXXXXXX : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX46, Y =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX16 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX0, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX2, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX21);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX2 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX3 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX2, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX4 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX3, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX5 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX4, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX5);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX6 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX5, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX6);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX7 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX6, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX7);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX8 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX7, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX8);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX9 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX8, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX9);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX10 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX9, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX10);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX11 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX10, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX11);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX12 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX11, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX12);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXXX13 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXXX12, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX13);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXX1 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXX8, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXXXXX : AXOI5 port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXXXXX1, C => XXXXXXXXXXXXXXXXXXXXXX
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXXXXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXX12 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX44, S => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXXXXXXX0, B
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX46);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX10 : AO1 port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXXXXX0, C => XXXXXXXXXXXXXXXXXXXXXX
                           , Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX20
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXX : NOR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXJXXXXXHXLXX, 
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXXXXXXXXXX : NOR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX0, Y
                           => XXXXXXXXXXXXXXXXXXXXXX5);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXX0 : NOR2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXX, Y =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXZXXXXXXXXXXXXX : OR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX0, B => XXXXXXXXXXXXXXXXXXXXXX
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXXXX : OR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP0, B =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXXXXXXX0 : OR3C port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXX2, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXX0 : OR3A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX11, 
                           B => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, C
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX1, 
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX15);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX : AO1B port map( A => 
                           MXMXXXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX1, C 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX, 
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX12);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX0 : AO1B port map( A => 
                           XXXXXXXX2, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX1, C 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX0,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX13);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX1 : OR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXX0, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX1,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXMXXX, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX14);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX2 : AO1B port map( A => 
                           MXMXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX1, C 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX2,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX16);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX3 : AO1B port map( A => 
                           MXMXXXXXXXX2, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX1, C 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX3,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX19);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXX1 : NOR3 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP0, C =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXX2 : NOR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX1, B
                           => XXXXXXXXXXXXXXXXXXXXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXXXXX : NOR3B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX0,
                           C => XXXXXXXXXXXXXXXXXJXXXXX1, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXJXXXXXHXLXXXXX : OR3C port map( A =>
                           XXXXXXXXXXXXXXXXXXXXXX5, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, C => 
                           XXXXXXXXXXXXXXXXXJXXX, Y => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX4 : AO1B port map( A => 
                           XXXXXXXX3, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2, C
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX4,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX15);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX5 : AO1B port map( A => 
                           XXXXXXXX4, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2, C
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX5,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX17);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX6 : AO1B port map( A => 
                           XXXXXXXX5, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2, C
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX6,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX18);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXX3 : NOR3 port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX0
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXX4 : NOR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX0, B => XXXXXXXXXXXXXXXXXXXXXX
                           , C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX3, Y
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX17 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX12, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX33)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX18 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX11, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX0
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX32);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX19 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX10, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX1
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX31);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX20 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX14, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX9, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX2
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX30);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX21 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX8, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX3
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX29);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX22 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX7, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX4
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX28);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX23 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX6, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX5
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX27);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX24 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX5, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX6
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX26);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX25 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX4, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX7
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX25);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX26 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX3, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX8
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX24);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX27 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX9
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX20);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXX28 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX16, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX29, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX10, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX7 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX9, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX7,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX11);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXX8 : AO1B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX8, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX8,
                           Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX10);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXX1 : OR3A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX12, 
                           B => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0
                           , C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2, Y
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX16);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXXXXXXX : NOR3B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX5, C => 
                           XXXXXXXXXXXXXXXXXJXXXXX2, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX0);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXXXX0 : NOR2A port map( A 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP0, B
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX4
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXXXX1 : NOR2A port map( A 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX4
                           , B => XXXXXXXXXXXXXXXXXXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXXXX2 : NOR2 port map( A =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX, B 
                           => XXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXXXXXXXXX : NOR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXP, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX3, 
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX11);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3 port map( A =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX3, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX, C
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX4, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX12);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX : AOI1B port map( A 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, B 
                           => XXXXXXXXXXXXXXXXXJXXXXX5, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX3, Y =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX9)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX0 : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX12, C 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX9,
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX6)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX1 : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX29, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0, 
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX, Y 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX10
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX2 : OA1A port map( A 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX35, C
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX10
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX5)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX3 : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX30, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0, 
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX0, Y
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX11
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX4 : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXXXX, C
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX11
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX4)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX5 : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0, B 
                           => XXXXXXXXXXXXXXXXXJXXXXX6, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXMXXX, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX12
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX6 : OA1A port map( A 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXX1, C
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX12
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX13
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX7 : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX4, 
                           B => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX13
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX14
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX8 : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX25, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0, 
                           C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX14
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX3)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX9 : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX7, C =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX15
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX2)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX10 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, B
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX8, C =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX16
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX0)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX11 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0, 
                           B => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX2, Y =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX17
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX12 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX26, 
                           B => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX0
                           , C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX17
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX18
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX13 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, B
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX9, C =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX18
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX : AOI1B port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXX0, Y 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX10);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX14 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX32, 
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX13,
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX19
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX15 : AOI1B port map( 
                           A => XXXXXXXXP0, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2, C
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX19
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX8)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX16 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX33, 
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX1, Y
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX20
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX17 : OA1A port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2
                           , B => XXXXXXXX1, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX20
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX7)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX0 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0, 
                           B => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXXXX44, C
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXXX, Y
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX9
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX1 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX36,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX3, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX8
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX2 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX37,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX4, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX7
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX3 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX38,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX5, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX6
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX4 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX39,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX6, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX5
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX5 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX40,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX7, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX4
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX6 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX41,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX8, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX3
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX7 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX42,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX9, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX2
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX8 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX43,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX10,
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX1
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX9 : AOI1B port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX44,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX11,
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX0
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXXX10 : AOI1B port map(
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX45,
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0,
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXX12,
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXX)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXXXXXXX : NOR3B port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX2, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX1, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, Y =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX : NOR3 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX2, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXXXX, C
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX3, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX2)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXXXXXXX0 : NOR3C port map( A =>
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX2, C 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXX0)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXXXXXXXXX : OR3 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX4, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX5, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX6, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXPXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX18 : NOR2A port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX2, B
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX21
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX19 : AND2 port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX0, B
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX21
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX1)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX20 : NOR2A port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX3, B
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX22
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX21 : AND2 port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX1, B
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX22
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX16
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX22 : NOR2A port map( 
                           A => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX4, B
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2, 
                           Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX23
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXXXXXXX23 : AND2 port map( A
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXMXXX, B 
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX23
                           , Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXVXXXXX15
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXX2 : NAND2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXX3 : NAND2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX1, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXXXXXXX4 : NAND2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXJXXXMXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXX7 : INV port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13, Y => 
                           XXXXXXXXXXXXXXXXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXXXX : OR3A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXXXX11, 
                           B => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, C
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2
                           , Y => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX14)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXX2 : OR3 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX2, B 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXX3, 
                           C => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX11, Y
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX17);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXX3 : OR2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX16);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXXXX4 : OR2 port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH, B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXH0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX15);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXXXXXXX : NOR3C port map( A 
                           => XXXXXXXXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXXXXXXXXXXXXXXXX, C => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX3, Y
                           => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX0)
                           ;
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX4, E => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXPXXX, CLK
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, CLR => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4, Q => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX13);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXHXLXXJXXXXX : BUFF port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX4);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXHXLXXJXXXXX0 : BUFF port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX3);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXHXLXXJXXXXX1 : BUFF port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX2);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXHXLXXJXXXXX2 : BUFF port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXX1);
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXXXX : NOR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXJXXXXXHXLXX, 
                           B => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX, Y 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXHXXXX2
                           );
   XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXHXLXXJXXXXXXX : BUFF port map( A => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXXX3);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX7 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX15);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX8 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX0, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX00);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX9 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX1, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX16);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX10 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX2, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX20);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX11 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX3, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX30);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX12 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX4, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX40);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX13 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX5, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX50);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX14 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX6, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXX0, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX60);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX7, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX23);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX8, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, CLK => XLX,
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX24);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX9, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, CLK => XLX,
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX25);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXX2 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX10, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, CLK => XLX,
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX26);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXX3 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX11, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, CLK => XLX,
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX27);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXX4 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX12, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, CLK => XLX,
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX28);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, CLK => XLX,
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX0, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, CLK => XLX,
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX0, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX1);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX1, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX2);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX2, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX6, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX3);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX4 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX3, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX7, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX4);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX5 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX4, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX7, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX5);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX6 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX5, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX7, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX6);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX7 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX6, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX7, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX7);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXX8 : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXJXXXXX7, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, CLK => XLX, 
                           CLR => XXXXXXXX7, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX8);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXPXWX : DFN1E1C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXXXXX4, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX0, CLK => XLX, 
                           CLR => XXXXXXXX7, Q => XXXXXPXWX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXPXXX : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXXXXX3, E => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, CLK => XLX, CLR => 
                           XXXXXXXX7, Q => XXXXXPXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXLXYXXXXX : DFN1E1C0 port map( D => 
                           XXXXXXXX1, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXYPXXXHXL, 
                           CLK => XLX, CLR => XXXXXXXX7, Q => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXLXY);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXYPX : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXL, CLK 
                           => XLX, CLR => XXXXXXXX7, Q => 
                           XXXXXXXXXXXXXXXXXXXXXXXXXYPX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXX, CLK
                           => XLX, CLR => XXXXXXXX7, Q => XXXXXXXX8);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXYPX0 : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXXXXXXX, E => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, CLK => XLX, CLR => 
                           XXXXXXXX7, Q => XXXXXXXXXXXXXXXXXXXXXXXXXYPX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXHXLXX, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXX0, 
                           CLK => XLX, CLR => XXXXXXXX, Q => XXXXXXXX00);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXP : DFN1E0C0 port map( D => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXPXXHXLXX, E => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX0, CLK => XLX, 
                           CLR => XXXXXXXX, Q => XXXXXXXXP0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3A port map( A => 
                           XXXXXXX0, B => XXXXXXXX1, C => XXXXXXXX00, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXPXXHXLXXXXV : AO1C port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, B => 
                           XXXXXXXXXXXXXXXXXXXXXX2, C => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXMXXX, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXPXXHXLXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXMXXXXXXXX : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, B => 
                           XXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXMXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXHXLXXXXXXX : OR2 port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX4, B => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXHXLXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXXXXX : AO1C port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, C => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXXHXL, Y =>
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXL);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXXHXLXXXXX : NOR2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX0, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXXHXL);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXXXXX : NOR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, B => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXXXXX : OR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX15, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX23, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX13);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX13, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXYPXXXHXLXXXXX : NOR2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXYPXXXHXL);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXXXXXXX : AO1C port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXX0, C => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXXHXL, Y =>
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXXXXXX0 : MX2A port map( A => 
                           XXXXXXX0, S => XXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXLXY, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX1 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX23, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX1, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX14);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX2 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX14, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX7, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX7);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXXXXX0 : NOR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXX0, B => XXXXXXXXXXXXXXXXXXXXXX5
                           , Y => XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXYPXXXHXLXXXXXXX : AO1A port map( A 
                           => XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXLXY, B => 
                           XXXXXXXX1, C => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXYPXXXHXLXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXXXXXXX0 : OR2B port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXXHXL, B =>
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXYPXXXHXLXX, 
                           Y => XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXXXXXXXXXXHXLXX
                           );
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXFLXXH : OA1A port map( A => XXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX, C => MXMPXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX3 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX15, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX4 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX16, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX1, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX1);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX5 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX17, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX2, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX2);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX6 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX18, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXX0, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX3);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX7 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX19, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX4, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX4);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX8 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX20, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX5, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX5);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX9 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX21, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX6, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX6);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX10 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX22, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX8, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX8);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX11 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX23, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX9, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX9);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX12 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX24, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX10, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX10);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX13 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX25, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX11, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX11);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX14 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX26, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXXX12, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX12);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXX : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX1, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX8, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX2, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX, B => 
                           XXXXXXXXXXXXXXXXXJXXXXX9, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX15 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX00, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX24, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX15);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX16 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX16, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX25, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX16);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX17 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX20, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX26, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX17);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX18 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX30, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX27, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX18);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX19 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX40, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX28, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX19);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX20 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX50, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX20);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX21 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX60, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX21);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX22 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX24, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX2, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX22);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX23 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX25, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX3, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX23);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX24 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX26, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX4, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX24);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX25 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX27, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX5, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX25);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXXX26 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX28, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX6, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXX26);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXX1 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX7, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX1);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXXXXXXX2 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX0, S => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXX8, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXXX2);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXXXXX0 : NOR3C port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX0, C => 
                           XXXXXXXXXXXXXXXXXJXXX, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXXXXXXX : NOR3 port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXXXXXX0, C => 
                           XXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX0);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXFLXXHXX : OA1A port map( A => XXXXXXX1, B =>
                           MXXXXXXXXXXXXXXXXXXXXXXX, C => MXMPXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXXXXXXX0 : OR2A port map( A => 
                           XXXXXXXXXXXXXXXXXXXXXXJXXXXXHXL, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXX0, Y => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXXJXXXXX);
   XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXXXXXXX : NOR2B port map( A => 
                           XXXXXXXXXXXXXXXXXJXXX0, B => XXXXXXXXXXXXXXXXXXXXXX5
                           , Y => XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXJXXXXX);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity XYXX0007 is

   port( XLXXPX, MXXXXXXXXXXXXXXXXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXXX0 : out 
         std_logic;  MXMXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXPXXXXXX, MXXXXXXXXXXXXXXXXXXFXXXHX : out std_logic
         ;  MXXXXXXXXXXXXXXXXXFXXXHXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXXXXX
         : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXYXLXXXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX0 :
         in std_logic;  MXXXXXXXXXXXXXXYXLXXXXXX0, MXXXXXXXXXXXXXXYXLXXXXXX1 : 
         out std_logic;  MXXXXXXXXXXXXXXXXPPMX, MXXXXXXXXXXXXXXXXXXMXMPXXXX : 
         in std_logic;  MXXXXXXXXXXXXXXYXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXXXXX7, 
         MXXXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXXXX9, 
         MXXXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXXXX11 : out std_logic
         ;  MXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXMWXXXXXXX, 
         MXXXXXXXXXXXXXXMWXXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXLLXX, 
         MXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXYXXXX, 
         MXXXXXXXXXXXXXXYXXXX0, MXXXXXXXXXXXXXXYXXXX1, MXXXXXXXXXXXXXXXXXFXXXHX
         , MXXXXXXXXXXXXXXYXLXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXPXXXXXX,
         MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, MXMXXXXXXXXXXXXXXX0, 
         MXMXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXMXMPXXXX, MXXXXXXXXXXXXXXXXXXXMXMPXXXX0, 
         MXXXXXXXXXXXXXXXXXXXPXXXXXX0, MXMXXXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXXXX3
         , MXXXXXXXXXXXXXMXMPXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0 : out std_logic;  
         MXMXXXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXXXX6, 
         MXMXXXXXXXXXXXXXXX7, MXMXXXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXXXPXXXXXX1, MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX9
         , MXXXXXXXXXXXXXXXXXXX0, XXXXXXXXXXXXXXXXXX : in std_logic;  MXVX : 
         out std_logic;  MXMXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX,
         MXMXXXXXXXXXXXXXXX11, MXMXXXXXXXXXXXXXXX12, MXMXXXXXXXXXXXXXXX13 : in 
         std_logic;  MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX : out std_logic;  
         MXMXXXXXXXXXXXXXXX14, MXMXXXXXXXXXXXXXXX15 : in std_logic;  
         MXXXXXXXXXXXXXXYXLXXXX0, MXXXXXXXXXXXXXXYXX : out std_logic;  
         MXMXXXXXXXXXXXXXXX16, MXMXXXXXXXXXXXXXXX17 : in std_logic;  
         MXXXXXXXXXXXXXXYXLXXXX1, MXXXXXXXXXXXXXXYXLXXXX2, MXXXXXXXXXXXXXXYXX0,
         MXXXXXXXXXXXXXXYXXXX2, MXXXXXXXXXXXXXXYXX1 : out std_logic;  
         MXMXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXMXMPXXXXXXX0, 
         MXXXXXXXXXXXXXMXMPXXXXXXX1 : in std_logic;  MXXXXXXXXXXXXXXXXYXLXXXXX 
         : out std_logic;  MXMXXXXXXXXXXXXXXX19, MXMXXXXXXXXXXXXXXX20, 
         MXXXXXXXXXXXXXXXXXXPXXLXX, MXXXXXXXXXXXXXXXXXMXVXWXXX, 
         MXXXXXXXXXXXXXXXXXXX1 : in std_logic;  MXXXXXXXXXXXXXXXXXXLL : out 
         std_logic;  XXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXPFF, MXMXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXX2, 
         MXMXXXXXXXXXXXXX3, MXMXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXX5, 
         MXMXXXXXXXXXXXXX6 : in std_logic;  MXXXXXXXXXXXXXXXXXX1 : out 
         std_logic;  MXXXXXXXXXXXXXMXMPXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXX : 
         in std_logic;  MXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXMWXXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX : in 
         std_logic;  MXXXXXXXXXXXXXXXXYXLXXXXX0, MXXXXXXXXXXXXXXXXYXLXXXXX1, 
         MXXXXXXXXXXXXXXXXYXLXXXXX2, MXXXXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXX2 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXX3 : in std_logic;  MXXXXXXXXXXXXXXXXXXXXX4, 
         MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXX6, 
         MXXXXXXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXXXXX8 : out std_logic);

end XYXX0007;

architecture SYN_USE_DEFA_ARCH_NAME of XYXX0007 is

signal MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXPXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXFXXXHX0, MXXXXXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX, MXXXXXXXXXXXXXXYXLXXXXXX2, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX0, MXXXXXXXXXXXXXXYXLXXXXXX00, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX1, MXXXXXXXXXXXXXXYXLXXXXXX10, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX, MXXXXXXXXXXXXXXXXPXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX
   , MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXXXX80, MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0, MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXX
   , MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX, MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXFXXXHX0, MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXMPXXX, 
   MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, MXXXXXXXXXXXXXXYXLXXXX3, 
   MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXMXVXXX, MXXXXXXXXXXXXXXXXPXXXXXXMXVXXX0, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXPXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXPXXXXXXX0, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX23, MXXXXXXXXXXXXXXXXPXXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXPXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXX0, MXXXXXXXXXXXXXXXXPXXXXXX1, 
   MXXXXXXXXXXXXXXXXPXXXXXX2, MXXXXXXXXXXXXXXXXPXXXXXX3, 
   MXXXXXXXXXXXXXXXXPXXXXXX4, MXXXXXXXXXXXXXXXXPXXXXXXX1, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXPXXXXXXX2, 
   MXXXXXXXXXXXXXXXXPXXXXXXX3, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXPXXXXXXX4, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXPXXXXXXX5, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXPXXXXXXX6, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXPXXXXXXX7, 
   MXXXXXXXXXXXXXXXXPXXXXXXX8, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXPXXXXXXX9, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXX1,
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXPXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXPXXXXXX5, 
   MXXXXXXXXXXXXXXXXPXXXXXX6, MXXXXXXXXXXXXXXXXPXXXXXX7, 
   MXXXXXXXXXXXXXXXXPXXXXXX8, MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX28, MXXXXXXXXXXXXXXXXPXXXXXX9, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX29, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXPXXXXXX10, 
   MXXXXXXXXXXXXXXXXPXXXXXX11, MXXXXXXXXXXXXXXXXPXXXXXXX10, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXPXXXXXX12, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXPXXXXXX13, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXPXXXXXXX11, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXX1, MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX16,
   MXXXXXXXXXXXXXXXXPXXXXXX14, MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXPXXXXXX15, MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXXPXXXXXX16, MXXXXXXXXXXXXXXXXPXXXXXXX12, 
   MXXXXXXXXXXXXXXXXPXXXXXXX13, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXPXXXXXXX14, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXPXXXXXXX15, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXXXPXXXXXXX16, 
   MXXXXXXXXXXXXXXXXPXXXXXXX17, MXXXXXXXXXXXXXXXXPXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXPXXXXXXX18, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXPXXXXXXX19, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXPXXXXXXX20, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXX, MXXXXXXXXXXXXXXXXPXXXXXXX21, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXX3, MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX00, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXXXXPXXXXXXX22, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX32, MXXXXXXXXXXXXXXXXPXXXXXXX23, 
   MXXXXXXXXXXXXXXXXPXXXXXXX24, MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXPXXXXXX17, MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXPXXXXXXX25, 
   MXXXXXXXXXXXXXXXXPXXXXXXX26, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXMXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX33, MXXXXXXXXXXXXXXXXPXXXXXXX27, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXPXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXPXXXXXX18, MXXXXXXXXXXXXXXXXPXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXX, MXXXXXXXXXXXXXXXXPXXXXXXX28, 
   MXXXXXXXXXXXXXXXXPXXXXXXX29, MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXPXXXXXXX30, 
   MXXXXXXXXXXXXXXXXPXXXXXXX31, MXXXXXXXXXXXXXXYXLXXXX00, MXXXXXXXXXXXXXXYXX2, 
   MXXXXXXXXXXXXXXXXPXXXXXXX32, MXXXXXXXXXXXXXXYXLXXXX10, 
   MXXXXXXXXXXXXXXXXPXXXXXXX33, MXXXXXXXXXXXXXXYXLXXXX20, 
   MXXXXXXXXXXXXXXXXYXLXXXXX3, MXXXXXXXXXXXXXXXXPXXXXXYXLXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXMXXX, MXXXXXXXXXXXXXXXXPXXXXXXXXM, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXX, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX, MXXXXXXXXXXXXXXXXPXXXXXXXM, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX0, MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX1, 
   MXXXXXXXXXXXXXXXXPXXXXXXXX2, MXXXXXXXXXXXXXXXXPXXXXXXMXMPXXXX, 
   MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX7, MXXXXXXXXXXXXXXXXPXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX2, MXXXXXXXXXXXXXXXXPXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXLL0, 
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXLLXXXXXXX, MXXXXXXXXXXXXXXXXYXLXXXXX00, 
   MXXXXXXXXXXXXXXXXYXLXXXXX10, MXXXXXXXXXXXXXXXXYXLXXXXX20, 
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXX, MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXX0, 
   MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX0, MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX1, 
   MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX2, MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX3, MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX4, MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX5, 
   MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX6, MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX7, 
   MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX0, MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX2 : std_logic;

begin
   
   MXXXXXXXXXXXXXXXXXXXPXXXXXX <= MXXXXXXXXXXXXXXXXXXXPXXXXXX2;
   MXXXXXXXXXXXXXXXXXXFXXXHX <= MXXXXXXXXXXXXXXXXXXFXXXHX0;
   MXXXXXXXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXXXXX0;
   MXXXXXXXXXXXXXXYXLXXXXXX <= MXXXXXXXXXXXXXXYXLXXXXXX2;
   MXXXXXXXXXXXXXXYXLXXXXXX0 <= MXXXXXXXXXXXXXXYXLXXXXXX00;
   MXXXXXXXXXXXXXXYXLXXXXXX1 <= MXXXXXXXXXXXXXXYXLXXXXXX10;
   MXXXXXXXXXXXXXXXXXXXXXXX8 <= MXXXXXXXXXXXXXXXXXXXXXXX80;
   MXXXXXXXXXXXXXXXXXFXXXHX <= MXXXXXXXXXXXXXXXXXFXXXHX0;
   MXXXXXXXXXXXXXXYXLXXXX <= MXXXXXXXXXXXXXXYXLXXXX3;
   MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX00;
   MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX <= 
      MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX0;
   MXXXXXXXXXXXXXXYXLXXXX0 <= MXXXXXXXXXXXXXXYXLXXXX00;
   MXXXXXXXXXXXXXXYXX <= MXXXXXXXXXXXXXXYXX2;
   MXXXXXXXXXXXXXXYXLXXXX1 <= MXXXXXXXXXXXXXXYXLXXXX10;
   MXXXXXXXXXXXXXXYXLXXXX2 <= MXXXXXXXXXXXXXXYXLXXXX20;
   MXXXXXXXXXXXXXXXXYXLXXXXX <= MXXXXXXXXXXXXXXXXYXLXXXXX3;
   MXXXXXXXXXXXXXXXXXXLL <= MXXXXXXXXXXXXXXXXXXLL0;
   MXXXXXXXXXXXXXXXXYXLXXXXX0 <= MXXXXXXXXXXXXXXXXYXLXXXXX00;
   MXXXXXXXXXXXXXXXXYXLXXXXX1 <= MXXXXXXXXXXXXXXXXYXLXXXXX10;
   MXXXXXXXXXXXXXXXXYXLXXXXX2 <= MXXXXXXXXXXXXXXXXYXLXXXXX20;
   
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXMXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX0, B => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXYXLXXXXXX : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX, CLK => XLXXPX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXYXLXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXYXLXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX0, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXYXLXXXXXX00);
   MXXXXXXXXXXXXXXXXPXXXYXLXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXYXLXXXXXX10);
   MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX, B => 
                           MXXXXXXXXXXXXXXXXPPMX, C => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX2, B => 
                           MXXXXXXXXXXXXXXYXLXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXYXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX7, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX4 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX5 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX6 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX80);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX7 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX8 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXX9 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX10, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXPXXXMWXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXMWXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXMWXXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXLLXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXX, E => MXXXXXXXXXXXXXXXXXXX, CLK 
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXLLXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX0, B => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX0, B => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX, B => 
                           MXXXXXXXXXXXXXXXXPPMX, C => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX2, B => 
                           MXXXXXXXXXXXXXXYXLXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX, Y => MXXXXXXXXXXXXXXYXXXX
                           );
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX2, B => 
                           MXXXXXXXXXXXXXXYXLXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXYXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX2, B => 
                           MXXXXXXXXXXXXXXYXLXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXYXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXFXXXHXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXFXXXHX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXLXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXMPXXX, B => 
                           MXXXXXXXXXXXXXXYXLXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXLXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, B 
                           => MXXXXXXXXXXXXXXYXLXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXFXXXHXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX3, B => 
                           MXXXXXXXXXXXXXXYXLXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXMXVXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXVXXX, B => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXVXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXMXVXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX80, B => 
                           MXXXXXXXXXXXXXXXXXFXXXHX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXVXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX0 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX3 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX4 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX1, B => MXMXXXXXXXXXXXXXXX0
                           , C => MXXXXXXXXXXXXXXXXPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX : OA1A port map( A => 
                           MXMXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX3 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX4 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXX4, S
                           => MXXXXXXXXXXXXXXXXPXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX25, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX5 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX6 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX0, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX7 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX28, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX8 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX10 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX1 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX2 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX5 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX6 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX7 : XAI1 port map( A => 
                           MXMXXXXXXXXXXXXXXX2, B => MXMXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX8 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX9 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX2, A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXX1, C 
                           => MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX19, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX0 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX00, B => 
                           MXMXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXXXXXXX : OR3 port map( A => 
                           MXMXXXXXXXXXXXXXXX4, B => MXMXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX0 : OR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX11 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX32);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX1 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX24, C => 
                           MXMXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXX : NOR3A port map( A => 
                           MXMXXXXXXXXXXXXXXX3, B => MXMXXXXXXXXXXXXXXX2, C => 
                           MXMXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX4, B => MXMXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX6, C => MXXXXXXXXXXXXXXXXPXXXXXXX9
                           , Y => MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX4 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX25, B => 
                           MXMXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX26, B => 
                           MXMXXXXXXXXXXXXXXX4, C => MXMXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX18, B => 
                           MXMXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX5 : NOR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX3, B => MXMXXXXXXXXXXXXXXXXX, Y =>
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX6 : NOR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX7, B => MXMXXXXXXXXXXXXXXXXX, C =>
                           MXXXXXXXXXXXXXXXXPXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXXXXXXX0 : OR3A port map( A => 
                           MXMXXXXXXXXXXXXXXX4, B => MXMXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXXXXXXX1 : OR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX4 : NOR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXMXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX33);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX12 : NOR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX31);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXXX : NOR3A port map( A => 
                           MXMXXXXXXXXXXXXXXX0, B => MXMXXXXXXXXXXXXXXXXX, C =>
                           MXMXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX7 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX21, B => 
                           MXMXXXXXXXXXXXXXXX3, C => MXMXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX8 : NOR2A port map( A => 
                           MXMXXXXXXXXXXXXXXXXX0, B => MXMXXXXXXXXXXXXXXX5, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXX1 : OR3 port map( A => 
                           MXMXXXXXXXXXXXXXXXXX0, B => MXMXXXXXXXXXXXXXXX2, C 
                           => MXXXXXXXXXXXXXXXXXXXPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXXXX9 : NOR3A port map( A => 
                           MXMXXXXXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXXXX2, C =>
                           MXMXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR2B port map( A =>
                           MXMXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXX1 : NOR2B port map( A => 
                           MXMXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, B => MXXXXXXXXXXXXXXXXPPMX
                           , C => MXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX5);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX19, C => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX4);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX00, C => 
                           MXMXXXXXXXXXXXXXXX1, Y => MXXXXXXXXXXXXXXXXPXXXXXX14
                           );
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX2 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX16);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX16);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXX, B => 
                           MXMXXXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX0 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX10, B => 
                           MXMXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX3 : OR3A port map( A => 
                           MXMXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX12);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX33, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX10);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX28, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX14);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX15);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX29);
   MXXXXXXXXXXXXXXXXPXXXXXXMXVX : NOR3B port map( A => MXXXXXXXXXXXXXXXXXXX0, B
                           => MXXXXXXXXXXXXXXXXPXXXXXXMXVXXX0, C => 
                           XXXXXXXXXXXXXXXXXX, Y => MXVX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX4 : OR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXPXXXXXX18
                           , C => MXXXXXXXXXXXXXXXXPXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX0 : OR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX5, C => MXMXXXXXXXXXXXXXXX5
                           , Y => MXXXXXXXXXXXXXXXXPXXXXXXX8);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX5 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX6 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX7 : OR3C port map( A => 
                           MXMXXXXXXXXXXXXXXX5, B => MXMXXXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX20);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX, B => 
                           MXXXXXXXXXXXXXXXXPPMX, C => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX11, B => MXMXXXXXXXXXXXXXXX8, Y =>
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX12, B => MXMXXXXXXXXXXXXXXX13, Y 
                           => MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX1 : OR3C port map( A => 
                           MXMXXXXXXXXXXXXXXX8, B => MXMXXXXXXXXXXXXXXX11, C =>
                           MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX8 : OR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX1, C => 
                           MXMXXXXXXXXXXXXXXX14, Y => MXXXXXXXXXXXXXXXXPXXXXXX9
                           );
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX9 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX00, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX13 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX10 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX13);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX11 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX22);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX2 : OR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXX1 : MX2B port map( A => 
                           MXMXXXXXXXXXXXXXXX13, S => MXMXXXXXXXXXXXXXXX8, B =>
                           MXMXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX17);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXMXXXX : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX12, S => MXMXXXXXXXXXXXXXXX8, B =>
                           MXMXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXMXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX12 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX27, B => 
                           MXMXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX15);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX13 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX5 : NOR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX27, C => 
                           MXMXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX00, B => 
                           MXXXXXXXXXXXXXXYXLXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX, Y => MXXXXXXXXXXXXXXYXX2)
                           ;
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX11 : NOR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX5);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX12 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX28);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX1 : OR3A port map( A => 
                           MXMXXXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXXXX16, C => 
                           MXMXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX19);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX6 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX14 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXX11);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX3, B => 
                           MXXXXXXXXXXXXXXYXLXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX33);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX10, B => 
                           MXXXXXXXXXXXXXXYXLXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX00, B => 
                           MXXXXXXXXXXXXXXYXLXXXX20, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXYXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXX1 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX00, B => 
                           MXXXXXXXXXXXXXXYXLXXXX20, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXYXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXX2 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX00, B => 
                           MXXXXXXXXXXXXXXYXLXXXX20, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX, Y => MXXXXXXXXXXXXXXYXX1)
                           ;
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXMXXXXXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXMXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXMXXXXXXXXXXXXXXX, C => MXXXXXXXXXXXXXMXMPXXXXXXX1,
                           Y => MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXX2 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXMXXXXXXXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXYXLXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXYXLXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXMXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXMXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXM);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXX1 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXX, A => 
                           MXXXXXXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXXXX19, Y =>
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXX2 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXX, A => 
                           MXXXXXXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXXXX20, Y =>
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXM, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXX0 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXM, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX3 : AO1D port map( A => 
                           MXMXXXXXXXXXXXXXXX20, B => MXMXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX17);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX4 : AO1D port map( A => 
                           MXMXXXXXXXXXXXXXXX20, B => MXMXXXXXXXXXXXXXXX19, C 
                           => MXMXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX32);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX15 : OR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX15, B => MXMXXXXXXXXXXXXXXX20, C 
                           => MXXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXMPXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, Y
                           => MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXMPXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX1 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXMPXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXX2 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXMPXXXX, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXMPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXMXMPXXXXXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXXXMXVXWXXX, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXMXMPXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXYXX2, B => MXXXXXXXXXXXXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXLLXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXLL0, B => MXXXXXXXXXXXXXXYXX2, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXLLXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXX4 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXMXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXFXXXHXX : OR2B port map( A => XXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXPFF, Y => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX16, B => MXMXXXXXXXXXXXXXXX19, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX14 : OR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX20, B => MXMXXXXXXXXXXXXXXX15, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXX10);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXX0 : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX11);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXMXXXXXXXXXXXXX0, B => MXMXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX9);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXX5 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX13);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX18, B => MXMXXXXXXXXXXXXXXX16, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX15 : NOR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX19, B => MXMXXXXXXXXXXXXXXX17, C 
                           => MXMXXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX21);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXX1 : OR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX19, B => MXMXXXXXXXXXXXXXXX16, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXX18);
   MXXXXXXXXXXXXXXXXPXXXXXXXMXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXXPXXXXXXXM
                           );
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX16 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX4, B => 
                           MXMXXXXXXXXXXXXXXX16, C => MXMXXXXXXXXXXXXXXX17, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX16 : NOR2A port map( A => 
                           MXMXXXXXXXXXXXXX0, B => MXMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX27);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX13 : AO1 port map( A => 
                           MXMXXXXXXXXXXXXX1, B => MXMXXXXXXXXXXXXX2, C => 
                           MXMXXXXXXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXXPXXXXXXX4)
                           ;
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXX : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX18, B => MXMXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX12);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX14 : OR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX16, B => MXMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX17 : OR2A port map( A => 
                           MXMXXXXXXXXXXXXX4, B => MXMXXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX24);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX18 : NOR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX18, B => MXMXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX25);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXXXXX3 : OR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX18, B => MXMXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX19 : OR2A port map( A => 
                           MXMXXXXXXXXXXXXX2, B => MXMXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX23);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX20 : NOR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX16, B => MXMXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX30);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXX7 : OR3B port map( A => 
                           MXMXXXXXXXXXXXXX4, B => MXXXXXXXXXXXXXXXXPXXXXXXX25,
                           C => MXMXXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXXXXXXXXXXX15 : AO1C port map( A => 
                           MXMXXXXXXXXXXXXX5, B => MXMXXXXXXXXXXXXX, C => 
                           MXMXXXXXXXXXXXXX0, Y => MXXXXXXXXXXXXXXXXPXXXXXXX26)
                           ;
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXX17 : AO1D port map( A => 
                           MXMXXXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXX3, C => 
                           MXMXXXXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXXPXXXXXX18);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXX2 : AXO1 port map( A => 
                           MXMXXXXXXXXXXXXX3, B => MXMXXXXXXXXXXXXX5, C => 
                           MXMXXXXXXXXXXXXX4, Y => MXXXXXXXXXXXXXXXXPXXXXXX8);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXX3 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX21, C => MXMXXXXXXXXXXXXX6,
                           Y => MXXXXXXXXXXXXXXXXPXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX0, B => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, Y => 
                           MXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXX5 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXMXXXXXXXXXXXXX0, C => MXXXXXXXXXXXXXMXMPXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXXXXXXXXXXX4 : NOR3A port map( A => 
                           MXMXXXXXXXXXXXXX1, B => MXMXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, B => 
                           MXXXXXXXXXXXXXXXXPPMX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXPPMXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXXXXXXXXXXXXXX21 : NOR2 port map( A => 
                           MXMXXXXXXXXXXXXX, B => MXXXXXXXXXXXXXXXXPXXXXXXXXX0,
                           Y => MXXXXXXXXXXXXXXXXPXXXXXXX31);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXLLXXXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXMWXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXMWXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXMWXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXLLXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXX, E => MXXXXXXXXXXXXXXXXXXX, CLK 
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXLL0);
   MXXXXXXXXXXXXXXXXPXXXYXLXXXX : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX, CLK => XLXXPX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXYXLXXXX00);
   MXXXXXXXXXXXXXXXXPXXXYXLXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX0, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXYXLXXXX10);
   MXXXXXXXXXXXXXXXXPXXXYXLXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXYXLXXXX3);
   MXXXXXXXXXXXXXXXXPXXXYXLXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXYXLXXXX20);
   MXXXXXXXXXXXXXXXXPXXXXXYXLXXXXX0 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, PRE => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX00);
   MXXXXXXXXXXXXXXXXPXXXXXYXLXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX0, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX10);
   MXXXXXXXXXXXXXXXXPXXXXXYXLXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXLXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX20);
   MXXXXXXXXXXXXXXXXPXXXXXYXLXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXYXLXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXX : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXX29, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, PRE => MXXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX7, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX4 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX5 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXX6 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX10, E => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXYXXXXXXXXXYX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXFXXXHXXXXXXXX : AOI1A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXFXXXHXXXXXXXX0 : AND2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXX0, B => 
                           MXXXXXXXXXXXXXXYXLXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXFXXXHXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXX0, B => 
                           MXXXXXXXXXXXXXXYXLXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXXXXXFXXXHXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXYXXXXXX, B => 
                           MXXXXXXXXXXXXXXYXLXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXXX : AOI1A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXXX0 : AOI1A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX20, B => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX5);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX3, B => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX4);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX3);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX3, B => 
                           MXXXXXXXXXXXXXXYXLXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX6);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX20, B => 
                           MXXXXXXXXXXXXXXYXLXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX4 : AOI1A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX5 : AND2A port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX10, B => 
                           MXXXXXXXXXXXXXXYXLXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX6 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX10, B => 
                           MXXXXXXXXXXXXXXYXLXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXXXXXX7 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX00, B => 
                           MXXXXXXXXXXXXXXYXLXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXLXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXLXXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX3, B => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXLXXXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXPXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXLXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX00, B => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXMPXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXLXXXXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX00, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX);
   MXXXXXXXXXXXXXXXXPXXXXXXXYXLXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX00, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXYXXLXXXXXXYXXX, Y => 
                           MXXXXXXXXXXXXXXXXPXXXWXXXXXXXXXXXXXXMPXXX);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity XYXX0006 is

   port( MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, XLXPXX, MXXXXXXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXFXWXXX, XFXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXPXWXXXXWXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXXX0 
         : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXXVXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXXX : out std_logic;  MXXXXXXXXXXXXXXXMXMXXXLXXXXXX
         , MXXXXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXXXX0 : out 
         std_logic;  MXXXXXXXXXXXXXXYXXXX, MXXXXXXXXXXXXXXYXXXX0 : in std_logic
         ;  MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9, MXXXXXXXXXXXXXXXXPXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12, MXXXXXXXXXXXXXXXXVXXXXXX, 
         MXXXXXXXXXXXXXXXXVXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXFX, 
         MXXXXXXXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXXXVXXXXXX1, 
         MXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXX0 : out std_logic;  
         MXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXL : out std_logic; 
         MXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXFX0 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXVXXXXXX2, 
         MXXXXXXXXXXXXXXXXVXXXXXX3, MXXXXXXXXXXXXXXXXXX1 : out std_logic;  
         MXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXX2 : in 
         std_logic;  MXXXXXXXXXXXXXXXXXXFXXXXX, MXXXXXXXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXXXPXXXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXFXWXXX : 
         in std_logic;  MXXXXXXXXXXXXXXXXXXX2 : out std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXXXPXXXXXXXX1, MXXXXXXXXXXXXXXXXPXXXXXXXX2 : out 
         std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX2, XXMXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXX4 : out std_logic;  XXXXX, MXXXXXXXXXXXXXXXXXXXXX2,
         XXXXX0, XXXX, XXXX0, XXXX1, XXXX2, XXXX3, XXXX4, 
         MXXXXXXXXXXXXXXXXXXXXX3 : in std_logic;  MXXXXXXXXXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXX4
         : out std_logic;  MXXXXXXXXXXXXXXXXXFXXXHXXX, MXXXXXXXXXXXXXXXXXFXXXHX
         , MXXXXXXXXXXXXXXFXXXXXXXXXXX1 : in std_logic;  XFXXXXXX : in 
         std_logic_vector (7 downto 0);  XFXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXXXXXXXX6 : in std_logic);

end XYXX0006;

architecture SYN_USE_DEFA_ARCH_NAME of XYXX0006 is

signal MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXWX, MXXXXXXXXXXXXXXXXXXXXXLXX, 
   MXXXXXXXXXXXXXXXXXXXXPXXXXXX0, MXXXXXXXXXXXXXXXXXXXLXXX0, 
   MXXXXXXXXXXXXXXXXXXXLXXX1, MXXXXXXXXXXXXXXXXXXXLXXXX, 
   MXXXXXXXXXXXXXXXXXXXLXXX2, MXXXXXXXXXXXXXXXXXXXLXXXXX, 
   MXXXXXXXXXXXXXXXXXXXLXXXXX0, MXXXXXXXXXXXXXXXXXXXLXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXLXXX3, MXXXXXXXXXXXXXXXXXXXX00, MXXXXXXXXXXXXXXXXXXXLX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX1, MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX2, MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX3, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX4, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, 
   MXXXXXXXXXXXXXXXXXXXXFXXPX, MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX6, 
   MXXXXXXXXXXXXXXXXXXXXXXXXPX, MXXXXXXXXXXXXXXXXXXXXFXXPX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXXXPX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXPX, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXXPX1, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX7, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXXPX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX8, MXXXXXXXXXXXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXX00, MXXXXXXXXXXXXXXXXXXXXXXXXLXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXX, MXXXXXXXXXXXXXXXXXXXXXXXXPXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX, MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXPXXX, MXXXXXXXXXXXXXXXXXXXXXXXPXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXLX, MXXXXXXXXXXXXXXXXXXXXXXXLXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX9, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXX1, MXXXXXXXXXXXXXXXXXXXXXXXXPXXX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXLXXX, MXXXXXXXXXXXXXXXXXXXXXXXXXPXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX1, MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX0, MXXXXXXXXXXXXXXXXXXXXXXXXPXXX2, 
   MXXXXXXXXXXXXXXXXXXXXFXXLX, MXXXXXXXXXXXXXXXXXXXXFXXPXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX1, MXXXXXXXXXXXXXXXXXXXXXXXLXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPX, MXXXXXXXXXXXXXXXXXXXXXXXPXXX1, 
   MXXXXXXXXXXXXXXXXXXXXFXXLX0, MXXXXXXXXXXXXXXXXXXXXFXXLXXX, 
   MXXXXXXXXXXXXXXXXXXXXFXXPXXX0, MXXXXXXXXXXXXXXXXXXXXXXXXLX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXX3, MXXXXXXXXXXXXXXXXXXXXXXXXPXXX4, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX10, MXXXXXXXXXXXXXXXXXXXXXXXXLXXX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX11, MXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, 
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXX6, MXXXXXXXXXXXXXXXXXXXXXXXXLX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXX3, MXXXXXXXXXXXXXXXXXXXLX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX2, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXXXXXLX3, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX4, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX5, MXXXXXXXXXXXXXXXXXXXXXXXXLX6, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX7, MXXXXXXXXXXXXXXXXXXXXXXXXXLX, 
   MXXXXXXXXXXXXXXXXXXXXPXXXX3, MXXXXXXXXXXXXXXXXXXXXFXXLX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXLX0, MXXXXXXXXXXXXXXXXXXXXXXXLX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX8, MXXXXXXXXXXXXXXXXXXXXFXXLX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXPXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX9, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX12, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX3, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX13, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX14, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX15, MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX0, 
   MXXXXXXXXXXXXXXXXXXXLX1, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX16, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXX4, MXXXXXXXXXXXXXXXXXXXXXXXXPXXX7, 
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXX8, MXXXXXXXXXXXXXXXXXXXXXXXXLX10, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX17, MXXXXXXXXXXXXXXXXXXXXXXXXLXXX5, 
   MXXXXXXXXXXXXXXXXXXXLXXX4, MXXXXXXXXXXXXXXXXXXXLXXX5, 
   MXXXXXXXXXXXXXXXXXXXLXXX6, MXXXXXXXXXXXXXXXXXXXLXXX7, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXX6, MXXXXXXXXXXXXXXXXXXXXXXXXLXXX7, 
   MXXXXXXXXXXXXXXXXXXXLXXXXX2, MXXXXXXXXXXXXXXXXXXXLXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXFXXLXXX0, MXXXXXXXXXXXXXXXXXXXLXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXXXXLXXX1, MXXXXXXXXXXXXXXXXXXXLXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXX8, MXXXXXXXXXXXXXXXXXXXXXXXXLXXX9, 
   MXXXXXXXXXXXXXXXXXXXXXXXLXXX2, MXXXXXXXXXXXXXXXXXXXXXXXXLXXX10, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX11, MXXXXXXXXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXLXXXXX6, MXXXXXXXXXXXXXXXXXXXLXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXLXXXXX8, MXXXXXXXXXXXXXXXXXXXXXXXXLX12, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXLX0, MXXXXXXXXXXXXXXXXXXXLXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXLXXXXX10, MXXXXXXXXXXXXXXXXXXXXXXXXLX13, 
   MXXXXXXXXXXXXXXXXXXXLXXXXX11, MXXXXXXXXXXXXXXXXXXXLXXXXX12, 
   MXXXXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXXPXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXXXXLX2, MXXXXXXXXXXXXXXXXXXXXXXXXLX14, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXPXXXX6, MXXXXXXXXXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXXXPXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXXXXPXXXX8, MXXXXXXXXXXXXXXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXPXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXXXXXXXXX21, MXXXXXXXXXXXXXXXXXXXLXXXXX13, 
   MXXXXXXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXX, 
   MXXXXXXXXXXXXXXXXVXXXXXX4, MXXXXXXXXXXXXXXXXVXXXXXX00, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXXXFF, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXFXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFF0, MXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFF1, MXXXXXXXXXXXXXXXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFF2, MXXXXXXXXXXXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXVXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXXXXXXPXXXX9, MXXXXXXXXXXXXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXX00, MXXXXXXXXXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFF3, MXXXXXXXXXXXXXXXXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFF4, MXXXXXXXXXXXXXXXL0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXXXXXXXXX27, MXXXXXXXXXXXXXXXXXXXXXXXX28, 
   MXXXXXXXXXXXXXXXXXXXXXXXX29, MXXXXXXXXXXXXXXXXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXXPX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXPX2, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXXXFXXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX5, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2, MXXXXXXXXXXXXXXXXXXXXXXXXPX3, 
   MXXXXXXXXXXXXXXXXXXXXXXXXPX4, MXXXXXXXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXVXXXXXX20, MXXXXXXXXXXXXXXXXVXXXXXX30, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX0, MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX1, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX2, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX18, 
   MXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFF5, MXXXXXXXXXXXXXXXXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFF6, MXXXXXXXXXXXXXXXXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXXXPXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX15, MXXXXXXXXXXXXXXXXXXXXXXXXLX16, 
   MXXXXXXXXXXXXXXXXXXXVXXXXXX1, MXXXXXXXXXXXXXXXXXXXXPXXXX11, 
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, MXXXXXXXXXXXXXXXXXXFXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXPXXXX12, MXXXXXXXXXXXXXXXXPXXXXXXXX00, 
   MXXXXXXXXXXXXXXXXXXXXPXXXX13, MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, 
   MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, MXXXXXXXXXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXXXXXXXLXXXXX14, 
   MXXXXXXXXXXXXXXXXXXXLXXXXX15, MXXXXXXXXXXXXXXXXXXXXXXXX32, 
   MXXXXXXXXXXXXXXXXXXXXXXXX33, MXXXXXXXXXXXXXXXXXXXVXXXXXXXX, 
   MXXXXXXXXXXXXXXXXPXXXXXXXX10, MXXXXXXXXXXXXXXXXPXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXXXXXXXXXLX17, MXXXXXXXXXXXXXXXXXXXXPXXXX14, 
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXVXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXVXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXXLX18 : std_logic;

begin
   MXXXXXXXXXXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXXXXXXX00;
   MXXXXXXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXXXX7;
   MXXXXXXXXXXXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXXXXXXXX00;
   MXXXXXXXXXXXXXXXXPXXXXXXXX <= MXXXXXXXXXXXXXXXXPXXXXXXXX3;
   MXXXXXXXXXXXXXXXXVXXXXXX <= MXXXXXXXXXXXXXXXXVXXXXXX4;
   MXXXXXXXXXXXXXXXXVXXXXXX0 <= MXXXXXXXXXXXXXXXXVXXXXXX00;
   MXXXXXXXXXXXXXXXXVXXXXXX1 <= MXXXXXXXXXXXXXXXXVXXXXXX10;
   MXXXXXXXXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXXXXX00;
   MXXXXXXXXXXXXXXXL <= MXXXXXXXXXXXXXXXL0;
   MXXXXXXXXXXXXXXXXXXXXX1 <= MXXXXXXXXXXXXXXXXXXXXX10;
   MXXXXXXXXXXXXXXXXVXXXXXX2 <= MXXXXXXXXXXXXXXXXVXXXXXX20;
   MXXXXXXXXXXXXXXXXVXXXXXX3 <= MXXXXXXXXXXXXXXXXVXXXXXX30;
   MXXXXXXXXXXXXXXXXXX1 <= MXXXXXXXXXXXXXXXXXX10;
   MXXXXXXXXXXXXXXXXXXFXXXXX <= MXXXXXXXXXXXXXXXXXXFXXXXX0;
   MXXXXXXXXXXXXXXXXPXXXXXXXX0 <= MXXXXXXXXXXXXXXXXPXXXXXXXX00;
   MXXXXXXXXXXXXXXXXXXX2 <= MXXXXXXXXXXXXXXXXXXX20;
   MXXXXXXXXXXXXXXXXPXXXXXXXX1 <= MXXXXXXXXXXXXXXXXPXXXXXXXX10;
   MXXXXXXXXXXXXXXXXPXXXXXXXX2 <= MXXXXXXXXXXXXXXXXPXXXXXXXX20;
   
   MXXXXXXXXXXXXXXXXXXXXPXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXLXX);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXXXXXFXWXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX, B => XFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX, C => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXPX, C => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX, C => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX, C => MXXXXXXXXXXXXXXXXXXXXX00,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX0 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX9, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXPXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX2);
   MXXXXXXXXXXXXXXXXXXXXFXXPXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXPX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPXXX1);
   MXXXXXXXXXXXXXXXXXXXXFXXPXXXXXXXX0 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX4 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX5 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX11, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX6 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX1, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX4 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX8, A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX7, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX12);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX5, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX13);
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX2, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX14);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX8, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX15);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX3, B => 
                           MXXXXXXXXXXXXXXXXXXXLX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX16);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX7 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX8);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX8 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX4 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX4, B => 
                           MXXXXXXXXXXXXXXXXXXXLX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX17);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX5 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX9, B => 
                           MXXXXXXXXXXXXXXXXXXXLX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX11);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX1, B => 
                           MXXXXXXXXXXXXXXXXXXXLX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX, B => MXXXXXXXXXXXXXXYXXXX0, C 
                           => MXXXXXXXXXXXXXXXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX6 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX10);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXX);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXX6);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXX1 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXX0);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXX1);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXX4);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXX4 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXX5);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXX5 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXX7);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX1);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX8, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX3);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX2 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX0);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX3 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX2);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX4);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX5);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX6 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX8);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX7 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLX0, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX10);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX8 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX13, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX1, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX12);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX7);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX6);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX11 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX9);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX12 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXVXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXX : NOR2B port map( A => MXXXXXXXXXXXXXXFX, 
                           B => MXXXXXXXXXXXXXXXXXXXXXLXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX16, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXLXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXLXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXX6 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXLX1);
   MXXXXXXXXXXXXXXXXXXXLXXX : OR3C port map( A => MXXXXXXXXXXXXXXXXXXXLXXXXX10,
                           B => MXXXXXXXXXXXXXXXXXXXLXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXLX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3C port map( A => MXXXXXXXXXXXXXXXXXX00
                           , B => MXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXLXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXLXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF4, B => 
                           MXXXXXXXXXXXXXXXL0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXX00, C => MXXXXXXXXXXXXXXXXXXX1
                           , Y => MXXXXXXXXXXXXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX27, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX);
   MXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX7 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX1);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXX : NOR3C port map( A => MXXXXXXXXXXXXXXXL0, B
                           => MXXXXXXXXXXXXXXFX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX8 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX9 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXLX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXVXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXVXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXVXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXVXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXLXXXXXX : OR3C port map( A => MXXXXXXXXXXXXXXXXXXXLXXX0,
                           B => MXXXXXXXXXXXXXXXXXXXLXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXLX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX15, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX1, B => 
                           MXXXXXXXXXXXXXXXXXXXLX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX);
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX0 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX3);
   MXXXXXXXXXXXXXXXXXXXXFXXPXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX1 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX2);
   MXXXXXXXXXXXXXXXXXXXXFXXPXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX2 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX17, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX10 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX11 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX18);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXX10, B => MXXXXXXXXXXXXXXXX0, C =>
                           MXXXXXXXXXXXXXXXL0, Y => MXXXXXXXXXXXXXXXXXXXXXXXXX0
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF5, B => 
                           MXXXXXXXXXXXXXXXL0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX4 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF6, B => 
                           MXXXXXXXXXXXXXXXL0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX3 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX13, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXPXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXPX);
   MXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLX0, B => MXXXXXXXXXXXXXXXXXXXLX
                           , Y => MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX9);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXPX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR2 port map( A => MXXXXXXXXXXXXXXXX1,
                           B => MXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXFXXLXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX);
   MXXXXXXXXXXXXXXXXXXXXFXXLXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX10);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX15);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX16);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX15, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX4 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX16, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX7);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX18, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX5 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXLXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX16, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX5);
   MXXXXXXXXXXXXXXXXXXXLXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXX00, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXL0, B => MXXXXXXXXXXXXXXXXXXFXXXXX0,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXXXXXFXWXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX00, B => MXXXXXXXXXXXXXXFXWXXX,
                           C => MXXXXXXXXXXXXXXXXXXFXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXWX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXXXXXFXWXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX00, B => MXXXXXXXXXXXXXXFXWXXX,
                           C => MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXFFXXXXXXXXXFXWXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX00, B => MXXXXXXXXXXXXXXFXWXXX,
                           C => MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXFFXXXXXXXXXFXWXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX00, B => MXXXXXXXXXXXXXXFXWXXX,
                           C => MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX1, B => MXXXXXXXXXXXXXXXXXXXXX00
                           , C => MXXXXXXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX1, B => MXXXXXXXXXXXXXXXXXXXXX00
                           , C => MXXXXXXXXXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX31);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX31, A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX28, B => 
                           MXXXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX32);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX1 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX1, B => MXXXXXXXXXXXXXXXXXXX0, Y
                           => MXXXXXXXXXXXXXXXXXXXXXXXX33);
   MXXXXXXXXXXXXXXXXXXXVXXXXXX : AOI1 port map( A => MXXXXXXXXXXXXXXXXXXXXXXXX3
                           , B => MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXXXXXFXWXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX6 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX9);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX4 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX9);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX7 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX5 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX1);
   MXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX12 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX6 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX2);
   MXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX8 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX17);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX9 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX2);
   MXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX0);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXXXX3 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXX3 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXFFXXXXXXXXFXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXXXXXFXXXXXXXXXXXXXXX : OR2A port map( A =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXFFXXXXXXXXFXXXXXXXXXXXXXXX0 : OR2B port map( A =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXXXXXFXXXXXXXXXXXXXXX0 : OR2 port map( A =>
                           XXMXXXXXXX, B => MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXFXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXXXX4 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXXXX5 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXX4 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXXXX6 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXX5 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXXX6 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX10 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX13);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX7 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX17, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX11 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX17, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX8);
   MXXXXXXXXXXXXXXXXXXXVXXXXXX0 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX1);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXX3 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXXPXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX0 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX18, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX13 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXPX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX14 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXFXXPX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX8);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXXXXX15 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXPX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX12 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX13 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX6);
   MXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX2 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXLX);
   MXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXPX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX8 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX18, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX8);
   MXXXXXXXXXXXXXXXXXXXXFXXLXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXFXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXPXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX14 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX7);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX15 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX12);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX9 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXLX);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX16 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX18, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX5);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX17 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX14);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXX);
   MXXXXXXXXXXXXXXXXXXXXFXXLXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXFXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX1);
   MXXXXXXXXXXXXXXXXXXXXFXXLXXXXXX2 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLX0);
   MXXXXXXXXXXXXXXXXXXXXFXXLXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXFXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXFXXLXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX18 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX11);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXX19 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLX18);
   MXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXX : DFN1C0 port map( D => XXXXX, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF4);
   MXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXX0 : DFN1C0 port map( D => XXXXX0, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF0);
   MXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXX1 : DFN1C0 port map( D => XXXX, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF5);
   MXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXX2 : DFN1C0 port map( D => XXXX0, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF3);
   MXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXX3 : DFN1C0 port map( D => XXXX1, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF);
   MXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXX4 : DFN1C0 port map( D => XXXX2, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF6);
   MXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXX5 : DFN1C0 port map( D => XXXX3, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF2);
   MXXXXXXXXXXXXXXXXXXXXXXXXFFXXXXX6 : DFN1C0 port map( D => XXXX4, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFF1);
   MXXXXXXXXXXXXXXXXXXXXXXXX0 : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, CLK => 
                           XLXPXX, PRE => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXX1 : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, CLK => 
                           XLXPXX, PRE => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX7, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX8, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX13 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXLX0, E => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX15);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX14 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXLX, E => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX13);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX15 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXLX1, E => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXXX3, Q => MXXXXXXXXXXXXXXXL0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXX0 : DFN1E1C0 port map( D => XFXXXXXX(0), E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXXX3, Q => MXXXXXXXXXXXXXXXXXX10)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX7 : DFN1E1C0 port map( D => XFXXXXXXXXXXX, E
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXXX3, Q => MXXXXXXXXXXXXXXXXXX00)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX8 : DFN1E1C0 port map( D => XFXXXXXX(3), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX9 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXVXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXVXXXXXX30);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXVXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXVXXXXXX00);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXX3 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXVXXXXXXXX0, E => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXVXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX32, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX33, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX29, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX33, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX33, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX30, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX33, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXXXXXPXXXX : DFN1E1C0 port map( D => XFXXXXXX(0), E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX : DFN1E1C0 port map( D => XFXXXXXXXXXXX, E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX11);
   MXXXXXXXXXXXXXXXXXXXXPXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX00);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX0 : DFN1E1C0 port map( D => XFXXXXXX(3), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX10);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX14);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX2 : DFN1E1C0 port map( D => XFXXXXXX(5), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX9);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX3 : DFN1E1C0 port map( D => XFXXXXXX(6), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX12);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX4 : DFN1E1C0 port map( D => XFXXXXXX(7), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX13);
   MXXXXXXXXXXXXXXXXXXXXPXXXX1 : DFN1E1C0 port map( D => XFXXXXXX(0), E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX5 : DFN1E1C0 port map( D => XFXXXXXX(1), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX8);
   MXXXXXXXXXXXXXXXXXXXXPXXXX2 : DFN1E1C0 port map( D => XFXXXXXX(2), E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX6 : DFN1E1C0 port map( D => XFXXXXXX(3), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX5);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX7 : DFN1E1C0 port map( D => XFXXXXXX(4), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX3);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX8 : DFN1E1C0 port map( D => XFXXXXXX(5), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX4);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX9 : DFN1E1C0 port map( D => XFXXXXXX(6), E =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX6);
   MXXXXXXXXXXXXXXXXXXXXPXXXXXXXXX10 : DFN1E1C0 port map( D => XFXXXXXX(7), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXXFXWX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXPXXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX10 : DFN1E1C0 port map( D => XFXXXXXX(0), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX11 : DFN1E1C0 port map( D => XFXXXXXX(1), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX12 : DFN1E1C0 port map( D => XFXXXXXX(2), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX13 : DFN1E1C0 port map( D => XFXXXXXX(3), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX14 : DFN1E1C0 port map( D => XFXXXXXX(4), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX15 : DFN1E1C0 port map( D => XFXXXXXX(5), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX16 : DFN1E1C0 port map( D => XFXXXXXX(6), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX17 : DFN1E1C0 port map( D => XFXXXXXX(7), E 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX2);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity XYXX0005 is

   port( MXXXXXXXXXXXXXXYXLXXXXXX, MXXXXXXXXXXXXXXYXLXXXXXX0 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXX1,
         MXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXX3 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXFXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0, 
         MXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1, MXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2
         : out std_logic;  MXXXXXXXXXXXXXXXXXXXFXWXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXFXWXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXFXWXXX
         , XFXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX0 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXFXWXXX0 : out std_logic;  XXXX : in std_logic;  
         MXXXXXXXXXXXXXXXX1 : out std_logic;  XXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX4 : in std_logic;  
         MXXXXXXXXXXXXXXXX2 : out std_logic;  MXXXXXXXXXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXYXLXXXXXX1, MXXXXXXXXXXXXXXYXLXXXX : in std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXMXXX : out std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
         XFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXX : 
         out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXWXXX, MXXXXXXXXXXXXXXLXXXVXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXFXWXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX3 : in std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXMXXX0 : out std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXXX, XFXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXXXXXXX7, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX8, MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX10, MXXXXXXXXXXXXXXFXXXXXXXXXXX11, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXXXXXXFXWXXX0 : in std_logic;  MXXXXXXXXXXXXXXXXXXMXXX, 
         MXXXXXXXXXXXXXXXXXXMXXXXX, MXXXXXXXXXXXXXXXXXXMXXX0 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXFXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXX1 : out std_logic;  XFXWX : in std_logic;  
         MXXXXXXXXXXXXXXFX : out std_logic;  MXXXXXXXXXXXXXXXXXXXX6 : in 
         std_logic;  MXXXXXXXXXXXXXXFX0 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXX7 : in std_logic;  MXXXXXXXXXXXXXXXXVXX : out 
         std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXPXWXXXXWXXX
         , XXMXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXMXXX1 : out std_logic
         ;  XXMXXXXXXX0, XXMXXXXXXX1, XLXPXX, MXXXXXXXXXXXXXXXXXXXXXXX, XX, XX0
         , MXXXXXXXXXXXXXXXXXXXXX : in std_logic;  XFXXXXXX : in 
         std_logic_vector (7 downto 1);  MXXXXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXX3 : in std_logic);

end XYXX0005;

architecture SYN_USE_DEFA_ARCH_NAME of XYXX0005 is

signal MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX1,
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX, MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, 
   MXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXX, MXXXXXXXXXXXXXXXXXMXXXXHXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX, MXXXXXXXXXXXXXXXXXMXXXXLXXXX,
   MXXXXXXXXXXXXXXXXXMXXXXLXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX3, MXXXXXXXXXXXXXXXXXMXXXXHXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, MXXXXXXXXXXXXXXXXXMXXXXLXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXXXFFX, MXXXXXXXXXXXXXXXXXMXXXXXXFFXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX1, MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX3, MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX5, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX6, MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXV1, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX0,
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX, MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX1, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX2
   , MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX3, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX4
   , MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX6, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX2, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX7, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX8
   , MXXXXXXXXXXXXXXXXXMXXXXLXXXX9, MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX10, MXXXXXXXXXXXXXXXXXMXXXXLXXXX10, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX4, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX11, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX12, MXXXXXXXXXXXXXXXXXMXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX5, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX13, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX14, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX6, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX16, MXXXXXXXXXXXXXXXXXMXXXXLXXXX11, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX7, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX18, MXXXXXXXXXXXXXXXXXMXXXXLXXXX12, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX8, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX19, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX20, MXXXXXXXXXXXXXXXXXMXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX9, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX21, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX22, MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX10, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX23, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX24, MXXXXXXXXXXXXXXXXXMXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX11, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX25, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX26, MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX12, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX27, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX28, MXXXXXXXXXXXXXXXXXMXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX13, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX29, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX30, MXXXXXXXXXXXXXXXXXMXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX14, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXV, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXX1, MXXXXXXXXXXXXXXXXXMXXXXHXXXX7, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX, MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX8, MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX2, MXXXXXXXXXXXXXXXXXMXXXXHXXXX9, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX10, MXXXXXXXXXXXXXXXXXMXXXXHXXXX11, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX3, MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX12, MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX6, MXXXXXXXXXXXXXXXXXMXXXXHXXXX13, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXX14, MXXXXXXXXXXXXXXXXXMXXXXLXXXLX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXX, MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX0, MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX3
   , MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX, MXXXXXXXXXXXXXXXXXMXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX5
   , MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX, MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX6, MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX0
   , MXXXXXXXXXXXXXXXXXMXXXXMXXXXX0, MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX7,
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX1, MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX8, MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX1
   , MXXXXXXXXXXXXXXXXXMXXXXXXXX1, MXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX1, MXXXXXXXXXXXXXXXXXMXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXX3, MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXX4, MXXXXXXXXXXXXXXXXXMXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX9, MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX1
   , MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX2, MXXXXXXXXXXXXXXXX00, 
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX3, MXXXXXXXXXXXXXXXXXMXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXX6, MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXX7, MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX11, 
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX12, MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX,
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX3, MXXXXXXXXXXXXXXXXXMXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX3, MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX13,
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX14, MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX0
   , MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX4, MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXXXFXWXXX2, MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX3, MXXXXXXXXXXXXXXXXXXFXWXXX00, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXX, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXXXX
   , MXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXXXX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX4,
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX5, MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX7, MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX8, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXX13, MXXXXXXXXXXXXXXXXXMXXXXLXXXX14, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX1, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX, MXXXXXXXXXXXXXXXXXMXXXXLXXXLX0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX2, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX0, MXXXXXXXXXXXXXXXXXMXXXXXXXPXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXMXXXXLXXXLXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX1, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX3, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX5, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX2, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX8, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX10, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX12, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXLXXXXXXX, MXXXXXXXXXXXXXXXXXMXXXXHXXXV, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX9, MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXV2, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX6, MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2, MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX10, MXXXXXXXXXXXXXXXXXMXXXXLXXXV, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLL, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX4, MXXXXXXXXXXXXXXXXXMXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXPXXXX, MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXLXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXLX, MXXXXXXXXXXXXXXXXXMXXXXHXXXV0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXX, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLL0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX1, MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXXXXXXFF0, MXXXXXXXXXXXXXXXXXMXXXXXXFFX0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXFXLL, MXXXXXXXXXXXXXXXXXMXXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX, MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFF, MXXXXXXXXXXXXXXXXXMXXXXXXXXFXLL, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFFX, 
   MXXXXXXXXXXXXXXXXXMXXXXLXXXVXFF, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLX0, MXXXXXXXXXXXXXXXXXMXXXXLXXXV0, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXFF, MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX1, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX2, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX3, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX4, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX5, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX7, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX8, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX9, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX10, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX11, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX12, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX28, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX13, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX29, 
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX14, MXXXXXXXXXXXXXXXXXMXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXX4, MXXXXXXXXXXXXXXXXXMXXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFF0, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFFX0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXLL0, MXXXXXXXXXXXXXXXXXMXXXXXXFXLL0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXFX1, MXXXXXXXXXXXXXXFX00
   , MXXXXXXXXXXXXXXXXXMXXXXHXXXVXFF0, MXXXXXXXXXXXXXXXXXMXXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX1, MXXXXXXXXXXXXXXXXXMXXXXLXXXVXFF0, 
   MXXXXXXXXXXXXXXXXXMXXXXXXFFXXXX, MXXXXXXXXXXXXXXXXXMXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXFXXXXXXXX, MXXXXXXXXXXXXXXXXXMXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXXXXXX0, MXXXXXXXXXXXXXXXXXMXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXXXXWXXXXFXXXXXXXXXX, MXXXXXXXXXXXXXXXXXMXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXXXXXXXX10 : std_logic;

begin
   MXXXXXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXXX8;
   MXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXX3;
   MXXXXXXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXXX00;
   MXXXXXXXXXXXXXXXXXXFXWXXX <= MXXXXXXXXXXXXXXXXXXFXWXXX2;
   MXXXXXXXXXXXXXXXXXXFXWXXX0 <= MXXXXXXXXXXXXXXXXXXFXWXXX00;
   MXXXXXXXXXXXXXXXX1 <= MXXXXXXXXXXXXXXXX10;
   MXXXXXXXXXXXXXXXX2 <= MXXXXXXXXXXXXXXXX20;
   MXXXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXX2;
   MXXXXXXXXXXXXXXFX <= MXXXXXXXXXXXXXXFX1;
   MXXXXXXXXXXXXXXFX0 <= MXXXXXXXXXXXXXXFX00;
   
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, C => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, C => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, C => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, C => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, C => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX2 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, C => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, C => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, B
                           => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX,
                           B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX
                           );
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0
                           , B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1
                           , B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, 
                           B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX,
                           Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, B
                           => MXXXXXXXXXXXXXXXXXMXXXXHXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, 
                           B => MXXXXXXXXXXXXXXXXXMXXXXHXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX5 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, 
                           B => MXXXXXXXXXXXXXXXXXMXXXXHXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0)
                           ;
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2
                           , B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2
                           );
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX,
                           B => MXXXXXXXXXXXXXXXXXMXXXXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX
                           , B => MXXXXXXXXXXXXXXXXXMXXXXLXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX5 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2
                           , B => MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX6 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3
                           , B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0
                           );
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX7 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX0, B =>
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3
                           );
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX8 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0
                           , B => MXXXXXXXXXXXXXXXXXMXXXXHXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX9 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXMXXXXHXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX10 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3
                           , B => MXXXXXXXXXXXXXXXXXMXXXXHXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX6 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4
                           , B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1
                           );
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX7 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX1, B =>
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4
                           );
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX8 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1
                           , B => MXXXXXXXXXXXXXXXXXMXXXXLXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX9 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, B 
                           => MXXXXXXXXXXXXXXXXXMXXXXLXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX10 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4
                           , B => MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXXXFFXXXXXXXX : INV port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXV : NAND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX6);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXX : NAND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXV1);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX,
                           C => MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX11 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX12 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX13 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX14 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX15 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX16 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX17 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX18 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX19 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX20);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX20 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX19);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX21 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX22);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX22 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX21);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX23 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX24);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX24 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX23);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX25 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX26);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX26 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX25);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX27 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX28);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX28 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX27);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX29 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX30);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXXXXXXX30 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX29);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXV, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX0);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX2);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX1);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXXXX3 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX4);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXXXX4 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX6);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXXXX5 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX5);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXXXX6 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX3 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX5 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX11);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX12);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX9 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX15);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX13);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX11 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX14);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXFFXXXXXXXXFXWXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXXXX0 : NOR2B port map( A => XFXXXXXXXXXX
                           , B => MXXXXXXXXXXXXXXFXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX00, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXXXXXXXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXX3, B => XXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXXXXXXXXX0 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXX10, B => XXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXXXX3 : NOR2B port map( A => XFXXXXXXXXXX
                           , B => MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXX3, B => MXXXXXXXXXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXX10, B => MXXXXXXXXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX5);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX7);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX8);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX1, B => 
                           MXXXXXXXXXXXXXXYXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXLXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXPXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX2 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX3 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX5 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, B => 
                           XFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX6 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX7 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX8 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX9 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX10 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX11 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX11);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX12 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, B => 
                           XFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX12);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX13 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX13);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXLXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX9);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXV2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX00, C => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXFFXXXXXXXXFXWX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXV0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX10);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXX : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLL, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXLX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXLXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXX3, C => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, Y => MXXXXXXXXXXXXXXXXXX2
                           );
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX00, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXLXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX4, B => 
                           MXXXXXXXXXXXXXXLXXXVXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXX0 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLL0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXX14 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX14);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXFXLLXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFF0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFXLL);
   MXXXXXXXXXXXXXXXXXMXXXXXXXPXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXPXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFF, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXLL, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLL0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXPXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXPXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFFXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFF, C => 
                           MXXXXXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFFX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXVXXXXX : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXV1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXVXFF, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXVXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXV2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXVXX10, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXXXXX1 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXFF, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXXXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX0, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX13);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX4 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX5 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX : MX2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX0 : MX2 port map( A => XFXXXXXXXXXXX0, S 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX5 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX6 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX6 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX7 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX14);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX8 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX11);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX9 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX10 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX11 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX12 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX12);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX13 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX7 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX8 : MX2 port map( A => XFXXXXXXXXXXX0, S 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX9 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX10 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX11 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX11);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX12 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX12);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX13 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX13);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXXXX14 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX14);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXLXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLXXX, B => 
                           MXXXXXXXXXXXXXXLXXXVXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXLXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXLXXXXX1 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXLXXXVXX, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFXLL, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXX : OR2B port map( A => MXXXXXXXXXXXXXXXX10, B
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXX : OR2B port map( A => MXXXXXXXXXXXXXXXX20,
                           B => MXXXXXXXXXXXXXXXXXMXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXLXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX12 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX13 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX14 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX15 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX16 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXFXXXXXXXMXXVXXXXXXXXXX17 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXFFXXXXXXXXFXWXXX0 : NOR2A port map( A => XFXWX
                           , B => MXXXXXXXXXXXXXXFXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXX3, B => MXXXXXXXXXXXXXXXXXXXX4, C 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLL, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFFXXXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFF0, C => 
                           MXXXXXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFFX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXXXXX0 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFF0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXLL0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLL);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXLXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXLXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFXLL0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXLX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX0 : MX2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX2 : MX2B port map( A => XFXXXXXXXXXXX0, S =>
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX3 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX6, B => 
                           MXXXXXXXXXXXXXXFX1, C => MXXXXXXXXXXXXXXXXXXXX6, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXFX00, C => MXXXXXXXXXXXXXXXXXXXX7, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXLXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXLX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXXXXXXX3 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXFF0, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXV : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV0, S => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXV, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV0, Y => 
                           MXXXXXXXXXXXXXXXXVXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXV, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXV, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXXXXXXX5 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXVXFF0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXFXLLXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFXLL0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXXXXXXX6 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXVXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXV);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXX10, B => MXXXXXXXXXXXXXXXXXXXX5, C 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLL0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFXLLXX0);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXFFXXXXXXXXFXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWXXXXXXXX3 : NOR2B port map( A => XFXWX, B => 
                           XXMXXXXXXX, Y => MXXXXXXXXXXXXXXXXXXFXWXXX00);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXX1 : OR2B port map( A => MXXXXXXXXXXXXXXFX00, 
                           B => MXXXXXXXXXXXXXXXXXMXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXXXXXXXXX0 : NOR2A port map( A => XXMXXXXXXX0
                           , B => XXMXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXFX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXXXX3 : OR3C port map( A => XXMXXXXXXX1, B 
                           => XXMXXXXXXX0, C => MXXXXXXXXXXXXXXXXXMXXXXLXXXX11,
                           Y => MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXLXXMXXXXXXXX3 : OR3C port map( A => XXMXXXXXXX1, B =>
                           XXMXXXXXXX0, C => MXXXXXXXXXXXXXXXXXMXXXXLXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXLXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXHXXMXXXXXXXX14 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXFXWX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXFFXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFX0, CLK => XLXPXX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFF0);
   MXXXXXXXXXXXXXXXXXMXXXXXXFFXXXXXX : DFN1C0 port map( D => XX, CLK => XLXPXX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXFF : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFXXX, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXFFXXXXXX0 : DFN1C0 port map( D => XX0, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXFFX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFFXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFF);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFFXXXXXX : DFN1C0 port map( D => XXXX0, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFFXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFF0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFFXXXXXX0 : DFN1C0 port map( D => XXXX, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFFX0);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXFFXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV0, E => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXFF0);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXVXFFXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXV, E => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXVXFF);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXVXFFXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV0, E => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXYXLX1, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXVXFF0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXVXFFXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXV, E => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXYXLX0, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXVXFF);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXLLXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFFX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXLL0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXFXLLXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXFFX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXLL);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX7, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX6, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX5, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX4, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX1 : DFN1E0C0 port map( D => XFXXXXXX(4), E
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX9, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXFX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXXXX3, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXXXX7, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXFX00);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXXXXX0 : DFN1E1C0 port map( D => XFXXXXXX(1), E
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXXXXX1 : DFN1E1C0 port map( D => XFXXXXXX(2), E
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXXXXX2 : DFN1E1C0 port map( D => XFXXXXXX(3), E
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXXXXX3 : DFN1E1C0 port map( D => XFXXXXXX(4), E
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXXXXX4 : DFN1E1C0 port map( D => XFXXXXXX(5), E
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXXXXX5 : DFN1E1C0 port map( D => XFXXXXXX(6), E
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXMXXXXXXXXXX6 : DFN1E1C0 port map( D => XFXXXXXX(7), E
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXFXWX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX7, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX8, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX9, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX10, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX11, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX12, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX13, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX14, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX13, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX12, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX11, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX10, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX13);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX14, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX9, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX8, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX7, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX12);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX9 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX1, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX10 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX2, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX13);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX11 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX3, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX12 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX4, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX11);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX13 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX5, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXHXXXXXXXXX14 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXXXX6, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX14);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX6, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX5, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX9 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX4, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX10 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX3, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX14);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX11 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX2, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX12 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX1, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX11);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX13 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX0, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXXXX14 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXXXXX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX12);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXFXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX0 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX1 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXFXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX3 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXX0 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXFXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX6 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXFXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX7 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXXX8 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXXLXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX11 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX12 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX13 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX14 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1
                           , Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX15 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX16 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX1, Y =>
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX17 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4
                           , Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX18 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX19 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX20 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX)
                           ;
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX11 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX12 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX13 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX14 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0
                           , Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX15 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX16 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX0, Y =>
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX17 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3
                           , Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX18 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX19 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX20 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXLXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXLXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX21 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX22 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX23 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX,
                           Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX25 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX
                           , Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX26 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX27 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2
                           , Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX28 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX29 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXXX30 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXLXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXLXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXMXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX21 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX22 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX23 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, Y
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX25 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, 
                           Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX26 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX27 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, 
                           Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX28 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2, Y 
                           => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX29 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0,
                           Y => MXXXXXXXXXXXXXXXXXMXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXXX30 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXXXXHXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXMXXXXXXXXHXXXLXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXXXXWXXXXXXXXXXXXXXMPXXX);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity XYXX0004 is

   port( XLXPXX, MXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX : in std_logic
         ;  MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXXXXXLXX, MXXXXXXXXXXXXXXLXXXVXX, 
         MXXXXXXXXXXXXXXXXXXXXX, XFXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX, 
         XFXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXLXXXXXXXXXX
         , MXXXXXXXXXXXXXXFXWXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX0 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXFXWXXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXXWXXX, MXXXXXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXX0 : out std_logic;  XFXXXXXXXXXX1, XXMXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXX, XFXXXXXXXXXXX, 
         XFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX5, MXXXXXXXXXXXXXXFXXXXXXXXXXX6, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX7, MXXXXXXXXXXXXXXFXXXXXXXXXXX8, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX9 : in std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXXX4 : out 
         std_logic;  MXXXXXXXXXXXXXXXXXXFXWXXX0, MXXXXXXXXXXXXXXXXXPXWXXXXWXXX,
         XFXWX, MXXXXXXXXXXXXXXXXVXX, XXMXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX1 
         : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXX6 : out std_logic;  MXXXXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXMXX, MXXXXXXXXXXXXXXLXXXVX, MXXXXXXXXXXXXXXLXXXVX0, 
         MXXXXXXXXXXXXXXXXXXXXXXXXX, XXXXX, MXXXXXXXXXXXXXXXXXXXXX0 : in 
         std_logic;  XXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX1 : in 
         std_logic;  XXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXX4, 
         MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXX6, 
         MXXXXXXXXXXXXXXXXXXXXX7 : in std_logic);

end XYXX0004;

architecture SYN_USE_DEFA_ARCH_NAME of XYXX0004 is

signal MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFFXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX,
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXLXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXX0, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX7,
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXX1, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX8,
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX11, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX14, MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXLXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX15, MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX16, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX17, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXLL, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXV, MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX0, MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXLXXX0, MXXXXXXXXXXXXXXXXXXFXWXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX18, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXLXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX20
   , MXXXXXXXXXXXXXXXXXXXXLXXXXXXX21, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX22, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX23, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX24, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX25, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX26, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX27, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX29, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX20, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX30, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX31, MXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX32, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX33, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34, MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXLXXXXXMP, 
   MXXXXXXXXXXXXXXXX00, MXXXXXXXXXXXXXXXXXXXXLXXXXXPXXXXMP, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXLXXXXXMP0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXPXXXXMP0, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX37, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX38, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX39, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX40, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX41, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX42, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX43, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXX, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX44, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX45, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX46, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX47, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX48, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX49, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX50, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXLL, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX51, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX15, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX23
   , MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX53, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMP, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXPXXXXMP, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXPXXXX, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXVXL, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXYXLX, MXXXXXXXXXXXXXXXXXXXXLXXXXXXYXLX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX54,
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX0, MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX2, MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX4, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX56, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX57, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX58, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFF, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXLXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFFXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXFFXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFF, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX0, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXX,
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX26,
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFXLL, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX28, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXMP, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX60, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX61, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX11, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX62, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX63, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX13, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX64, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX14, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX65, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX15, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX67, MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX68, MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX69, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX29, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX31, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX70, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX71, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX72, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX73, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX74, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX32, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX75, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXXLXXXXVXFF
   , MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXVXX, MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX6, MXXXXXXXXXXXXXXXXXXXXLXXXXXXXYXLX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMPXXXX, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX77, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXMPXX, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX79, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX80, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXLX, MXXXXXXXXXXXXXXXXXXXXLXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX81, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXX82, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX34, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXXXLXXXXXXX83, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4 : std_logic;

begin
   
   MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX0;
   MXXXXXXXXXXXXXXXXXXFXWXXX <= MXXXXXXXXXXXXXXXXXXFXWXXX1;
   MXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXX1;
   MXXXXXXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXXX00;
   
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX4, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXX, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX, CLK => XLXPXX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX
                           , B => MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXX,
                           Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX11, C
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX, B =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX, 
                           B => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX
                           );
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX
                           , B => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX8, Y =>
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFFXXXXXXX : INV port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFFXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX : AO1D port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX0 : AO1D port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX1 : AO1D port map( A 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX4, B 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3A port map( A
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3B port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3B port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXX : NOR3A port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX3
                           );
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXLXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXLXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3 port map( A
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX4
                           );
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXLXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXX1, B =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXXXX : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXXXX1, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX4)
                           ;
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3C port map( 
                           A => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX11, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3A port map(
                           A => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX : OA1 port map(
                           A => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXLXXXVXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXXXXXXXX : NOR2B port map( 
                           A => MXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXXX
                           );
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX3, B =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX4, Y =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX6, Y =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXXXX0 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXXXXXX : NOR3A port map( A => 
                           XFXXXXXXXXXX, B => MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           XFXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVX, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXXXX1 : NOR3C port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXLL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXXXXXXX : OR2 port map( A 
                           => MXXXXXXXXXXXXXXLXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXX0
                           );
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXXXXXXXXX : NOR2B port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXV, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXWXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR2 port map( 
                           A => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXLX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXLXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXLXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX18);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX11, C
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXLXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXLXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX, Y
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX22);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX1, 
                           Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX25);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX4
                           , C => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX26);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXXX
                           , B => MXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX27);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXX4, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX1 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXX0, 
                           A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX4, B 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX29);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX30);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXFXLLXXXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX33);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX7, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX0 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX5, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX1 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX6, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX2 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX3 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMP, B => 
                           MXXXXXXXXXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXPXXXXMP, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX1 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMP0, B => 
                           MXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXPXXXXMP0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX12, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6,
                           Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXLXXXXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX38, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX4, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXX2, B =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3B port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX41, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX5, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX42);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX43, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX40);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX44, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX32, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX45);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX46, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX47, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX48);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXX0 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX49, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX6, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX38);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX26, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX50, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXLL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX51, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX4, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX5, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXX2 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX50);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXX2 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX16);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX43, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX2 : OR2A port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX3 : OR2 port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX5, A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXXXX : NOR2A port map( A => XFXXXXXXXXXX1
                           , B => XXMXXXXXXX, Y => MXXXXXXXXXXXXXXXXXXFXWXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX9, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX9, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX4 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX9, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX53);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXPXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMP, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXPXXXXMP, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXPXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX24, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXPXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXVXL, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXYXLXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMP0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXYXLX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXYXLXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMP, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXYXLX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX : MX2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52, B => XFXXXXXXXXXXX,
                           Y => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX0 : MX2C port map( A => 
                           XFXXXXXXXXXXX0, S => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52
                           , B => MXXXXXXXXXXXXXXFXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX3 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX54, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX25, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXMXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXMXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX2 : MX2B port map( A => XFXXXXXXXXXXX0, S 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX0, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX1, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX2, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX3, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXXXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX4, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX56, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXLXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXLXXXXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX57, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX58);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFF, B => 
                           MXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX5 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX24);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX6 : NOR2 port map( A => 
                           XFXXXXXXXXXXX0, B => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34
                           , Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX23);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX7 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX21);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXXXXXX8 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXLXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX56, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXLXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXFFXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFFXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXFFXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFF, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFF, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX51);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX34);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXX : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXX0
                           , B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXX, C
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXFXLLXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFXLL, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXXXX, S
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLXXXXXXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX28, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXVXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0, S 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX54);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXX2 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX53, A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX30, A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXMP, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX60);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX61);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX62);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX63);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX13, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX64);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX14, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX65);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX15, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX67);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXXX5 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX16, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX68);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXXX6 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX17, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX69);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXLL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXLL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX4 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXLL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXLL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX31, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX70, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX71, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX37);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXX0 : OR2B port map( A => XFXWX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX55);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX43);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXLXXXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFXLL, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX32);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXFXLLXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX31);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXLXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX72, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX26, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX70);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX73, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX74, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX1 : NOR3B port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX73, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OR3B port map( A
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX75, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX10, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX50, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX2 : NOR3B port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX3 : NOR3A port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXV : NOR2A port map( A => MXXXXXXXXXXXXXXXXVXX,
                           B => MXXXXXXXXXXXXXXXXXXXXLXXXXVXFF, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXVXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX1 : NOR2B port map( A => 
                           XXMXXXXXXX0, B => MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXXXXXX5 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX5, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXFXXXXXXXXXXXX6 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXYXLXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMP, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXYXLX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMPXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX57, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMP, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMPXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXMPXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX45, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX77, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMPXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX47);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX79, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX80);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX49, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX79);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX80, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX44, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX71);
   MXXXXXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXMXXXXX, Y =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX41);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX43, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX17);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX44);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX42, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX38, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX49);
   MXXXXXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXMXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXLX, S => 
                           MXXXXXXXXXXXXXXMXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66);
   MXXXXXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXMX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXLXXXVX, S => MXXXXXXXXXXXXXXMXX, B =>
                           MXXXXXXXXXXXXXXLXXXVX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX81);
   MXXXXXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX81, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXMXXXXX, Y =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX72);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXFXWXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX52);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXLXXXXXXMX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXLXXXVX0, S => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX56);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVX, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX72, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX39);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXMXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX57);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXMXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX57, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX77);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX46);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX4 : NOR3B port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX74, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX5 : NOR3C port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX74, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3A port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX82, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXX1 : NOR3A port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX75, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR3B port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX82, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXX3 : NOR3B port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX75, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXX1 : NOR3C port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX76);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR3B port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX73);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OR2B port map( 
                           A => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX34, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX75);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR2 port map( A
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX34, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX74);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXX3 : OR2A port map( A 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX32);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : OR2A port map( 
                           A => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX34, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX82);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX82, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX9, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX6 : NOR3A port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX73, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX75, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX7 : NOR3A port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX73, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXX3, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXX8 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXXXX3, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXX1 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX82, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXXXXX4, C 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX5
                           );
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX74, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX3
                           , C => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX1 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX3, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX5, C
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXXXX3 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX51, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXXXXXXXXXXXXXXXX4 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX, S 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXX66, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX83);
   MXXXXXXXXXXXXXXXXXXXXLXXXXVXFFXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXVXX, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXVXFF);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFFXXXXX : DFN1P0 port map( D => XXXXX, CLK => 
                           XLXPXX, PRE => MXXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFFXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXX1, CLK => XLXPXX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFF);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFF : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFFXX, CLK => XLXPXX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFFXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXVXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXVXX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXLLXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXFFXXXXXXXXXXXX, 
                           CLK => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXLL);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX5, CLK
                           => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFXLLXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX6, CLK
                           => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFXLL);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXLLXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX4, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXLL);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXLXXXXXXXXXX, CLK
                           => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXLX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0, CLK => 
                           XLXPXX, PRE => MXXXXXXXXXXXXXXXXXXXXX0, Q => XXXXX0)
                           ;
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXVXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXLXXXXXXXXXX0, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXV);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXMPXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXLXXX0, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMP);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXMPXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMPXX, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMP0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFFXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXFF);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX32, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX58, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXX, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX48, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXFXLLXX, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX, CLK => XLXPXX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXPXXXXMPXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMP0, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXYXLX, CLK => XLXPXX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXPXXXXMP0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXPXXXXMPXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXMP, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXYXLX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXPXXXXMP);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXLXXXXX : DFN1E0P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX18, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXX, CLK => 
                           XLXPXX, PRE => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX : DFN1E0P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX83, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX14, CLK => 
                           XLXPXX, PRE => MXXXXXXXXXXXXXXXXXXXXX1, Q => XXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXPXXXXMPXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMP, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXYXLX, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXPXXXXMP);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX19, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXFXWX0, CLK => XLXPXX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXVXLXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXL, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX57, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXVXL);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMPXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMPXXXX, CLK => XLXPXX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXMP);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXMPXXXXX : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX27, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXMP);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX1, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX0 : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX27, CLK =>
                           XLXPXX, PRE => MXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX26, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX19, CLK =>
                           XLXPXX, PRE => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX20, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX23, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX22, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX24, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX21, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXXXXXXXX5
                           , CLK => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX25, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX10, CLK 
                           => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX5, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX6, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX7, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX8, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX9, CLK =>
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX0 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX11, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX1 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX12, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX2 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX13, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX3 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX14, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX4 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX15, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX5 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX16, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX6 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX17, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX7 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX60, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX78, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX17);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX8 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXX5, E =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX9 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX10 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX11 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX25, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX12 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX7, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX13 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX22, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX14 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX15 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX16 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX29, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXX17 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXX4 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXVXXXX, E =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX28, CLK => XLXPXX, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX61, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX4, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX62, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX63, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX64, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX65, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXX4 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX67, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXX5 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX68, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXXXXXXX6 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX69, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXX59, CLK => XLXPXX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXFXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXX : DFN1E0P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, CLK => XLXPXX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXX0 : DFN1E0P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, CLK => XLXPXX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXX1 : DFN1E0P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, CLK => XLXPXX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX9 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX4, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX10 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX5, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX11 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXXX5, CLK 
                           => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXXXXX12 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXXXX6, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1, 
                           CLK => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX5, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX6, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX7, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX7, CLK
                           => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX8, CLK
                           => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX9, CLK
                           => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX10, 
                           CLK => XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX11, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX12, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX13, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX13, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX14, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX15, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX16, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX9 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX4, CLK => 
                           XLXPXX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX2 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, C 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX3 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX
                           , B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX1, C 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX6 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX1, 
                           Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX7 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX8 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX9 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXXX10 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXX : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX
                           );
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXX0 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHXFXXXXXXXXXXXXX3 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXHXFXXXLX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX
                           , Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX31);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX29);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX4 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX, 
                           Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX,
                           Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX, Y =>
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX6 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, C 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX1 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXX, C 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX34);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX
                           , B => MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXX,
                           Y => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX33);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX8, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX6 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y =>
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX7 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX
                           );
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXX8 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX7, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX7, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX4 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX5 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX7, B 
                           => MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y
                           => 
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXX6 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXVXLXXXXXXXX0, Y =>
                           MXXXXXXXXXXXXXXXXXXXXLXXWXXXXXXXXXXXXXXMPXXX);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity XYXX0003 is

   port( MXXXXXXXXXXXXXXXXXXXXXX, XLXXPX, MXXXXXXXXXXXXXXXXXXXXXXXXX : in 
         std_logic;  XFXXXXXXXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX : 
         in std_logic;  XFXXXXXXXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXMXMPXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXPXXXXXX : out 
         std_logic;  MXXXXXXXXXXXXXXXXXXXPXXXXXX0 : in std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXXXXX : out std_logic;  MXMXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX : out std_logic;  MXMXXXXXXXXXXXXX0 
         : in std_logic;  MXXXXXXXXXXXXXXXXXXXPXXXXXX1 : out std_logic;  
         MXXXXXXXXXXXXXMXMPXXXXXXX, MXMXXXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXXXX0
         , MXMXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXX1, 
         MXMXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXX,
         MXXXXXXXXXXXXXXFXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXX5, 
         XFXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX6, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX7, XFXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX8, MXXXXXXXXXXXXXXFXXXXXXXXXX9, 
         XFXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXX0 : out std_logic;  
         MXXXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX2 : out std_logic;  MXXXXXXXXXXXXXXXXXX0 : 
         in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX4 : out std_logic;  MXXXXXXXXXXXXXXXXXX1 : 
         in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX6 : out std_logic;  MXXXXXXXXXXXXXXXXXX2 : 
         in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX7, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX8 : out std_logic;  MXXXXXXXXXXXXXXXXXX3 : 
         in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX10 : out std_logic;  MXXXXXXXXXXXXXXXXXX4 :
         in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX11 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXXX1 : in std_logic;  MXXXXXXXXXXXXXXFXWXXX : out
         std_logic;  MXXXXXXXXXXXXXXXXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX : out std_logic;  
         MXMXXXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXXXXXXXXXX3, XXXXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXPXXXXXXXX, XXXXXXX, XFXXXXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXYXXXX, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, 
         MXMXXXXXXXXXXXXXXX3, XFXXXXXXXXXXX, MXMXXXXXXXXXXXXXXX4, 
         MXXXXXXXXXXXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX6, 
         MXXXXXXXXXXXXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXXXX7, MXMXXXXXXXXXXXXXXX8, 
         MXMXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXMXMPXXXXXXX0 : in std_logic;  
         MXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXMXMPXXXX, 
         MXXXXXXXXXXXXXXXXXXXMXMPXXXX0, MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX : out 
         std_logic;  MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXPXXXX : out std_logic;  MXMXXXXXXXXXXXXXXX10 : in 
         std_logic;  MXXXXXXXXXXXXXXXXXX6 : out std_logic;  XXMXXXXX : in 
         std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0 : in std_logic;
         MXXXXXXXXXXXXXXXXXX7 : out std_logic;  XXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXX8 : out std_logic;  XXXXXXXX0 : in std_logic;  
         MXXXXXXXXXXXXXXXXXX9 : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX0 : in 
         std_logic;  MXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXX11, 
         MXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXX13 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  XXMXXXX
         : out std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXXYXXXX0, 
         MXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXVXXXXXX, XXXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXXXX2, XXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXVXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXXXVXX, MXXXXXXXXXXXXXXXXXXXXXXXVXX0, 
         MXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXX5 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXPXXXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX6
         , MXXXXXXXXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXXXXXXX8 : in std_logic;
         MXXXXXXXXXXXXXXXXXX14 : out std_logic;  MXXXXXXXXXXXXXXXXXX15, 
         MXXXXXXXXXXXXXXXXXXFXWXXX, MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, 
         MXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXXXX11 :
         in std_logic;  MXXXXXXXXXXXXXXXXXXFXXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXXWXXX, MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0, 
         XXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXFXWXXX0 : 
         in std_logic;  XFXXXXXX : out std_logic_vector (7 downto 2);  
         MXXXXXXXXXXXXXPXHXXXXXX : in std_logic;  XXMXXXXX0 : out 
         std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXPXHXXXXXX0, 
         MXXXXXXXXXXXXXPXHXXXXXX1, MXXXXXXXXXXXXXPXHXXXXXX2, 
         MXXXXXXXXXXXXXPXHXXXXXX3, MXXXXXXXXXXXXXPXHXXXXXX4, 
         MXXXXXXXXXXXXXPXHXXXXXX5, MXXXXXXXXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXFXWXXX1, 
         MXXXXXXXXXXXXXPXHXXXXXX6, MXXXXXXXXXXXXXXXXXXFXWXXX2, 
         MXXXXXXXXXXXXXMXMPXXXXXXX1, MXXXXXXXXXXXXXXYXXXX1, 
         MXXXXXXXXXXXXXXXXXXX6, XXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX1 : in
         std_logic;  MXXXXXXXXXXXXXXXXXXX7 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  XFXXXXXXXXXXXXXXXXX, 
         XFXXXXXXXXXXXXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXXXXXX9, 
         MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXMXMXMXXXX, 
         MXMXXXXXXXXXXXXXXX12, MXMXXXXXXXXXXXXXXX13, MXMXXXXXXXXXXXXXXX14, 
         MXMXXXXXXXXXXXXXXX15 : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXX : out 
         std_logic;  MXXXXXXXXXXXXXXXMXXX, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX, 
         MXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX,
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0, MXXXXXXXXXXXXXXXXXX17, 
         MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX, MXXXXXXXXXXXXXXXMXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1
         , MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2, 
         MXXXXXXXXXXXXXXXXXXMXXX, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXX, MXXXXXXXXXXXXXPXLXXXXXX, 
         MXXXXXXXXXXXXXPXLXXXXXX0, MXXXXXXXXXXXXXPXLXXXXXX1, 
         MXXXXXXXXXXXXXPXLXXXXXX2, MXXXXXXXXXXXXXPXLXXXXXX3, 
         MXXXXXXXXXXXXXPXLXXXXXX4, MXXXXXXXXXXXXXPXLXXXXXX5, 
         MXXXXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXX9, 
         MXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX0, MXXXXXXXXXXXXXXYXXXXXX, 
         MXXXXXXXXXXXXXXXXXXX10 : in std_logic;  XXMXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXX7, 
         MXMXXXXXXXXXXXXXXX16, MXMXXXXXXXXXXXXXXX17, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXX2, MXXXXXXXXXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXPXXXXXXX : in std_logic;  XFXXXXXX0 : in 
         std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXMXXX, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXPXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXPXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXPXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXX, MXXXXXXXXXXXXXXFXXXXXPXXXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXX4, XFXXXXXXXXXXX0, MXXXXXXXXXXXXXXXMXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1, MXXXXXXXXXXXXXXXXXX19, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3, MXXXXXXXXXXXXXXXXXX20, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXX2, MXXXXXXXXXXXXXXXMXXX2, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2, MXXXXXXXXXXXXXXXXXXX11, 
         MXXXXXXXXXXXXXXYXXXX2, MXXXXXXXXXXXXXXYXX, MXXXXXXXXXXXXXXXXXXX12, 
         MXXXXXXXXXXXXXMXMPXXXXXXX2, MXXXXXXXXXXXXXXXXXXMXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8, MXXXXXXXXXXXXXPXLXXXXXX6, 
         MXXXXXXXXXXXXXXXXXX21, MXMXXXXXXXXXXXXXXX18, MXMXXXXXXXXXXXXXXX19 : in
         std_logic;  MXXXXXXXXXXXXXXXXXX22, XFXWX : out std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5, MXXXXXXXXXXXXXXFXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXX3, MXXXXXXXXXXXXXXFXXXXXXXMXXX0, 
         MXXXXXXXXXXXXXXXXXX23, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10,
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7, MXXXXXXXXXXXXXXXMXXX3, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3, MXXXXXXXXXXXXXXXXXXMXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8
         , MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9, MXXXXXXXXXXXXXXXXXXXHXXX, 
         MXXXXXXXXXXXXXXXXXXFXWX, MXXXXXXXXXXXXXXXMXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4, MXXXXXXXXXXXXXXXXXXMXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11, MXXXXXXXXXXXXXXXXXXXHXXX0, 
         MXXXXXXXXXXXXXXXMXXX5, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2, MXXXXXXXXXXXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXX3, MXMXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12, MXXXXXXXXXXXXXXXXXX24, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12, MXXXXXXXXXXXXXXFXXXXXXLXXXX4, 
         MXXXXXXXXXXXXXXXMXXX6, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXX4, MXMXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXX5, 
         MXMXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXYXX0, MXXXXXXXXXXXXXXXXXX25, 
         MXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXX9 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXPXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX10
         , MXXXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXX26, 
         MXXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXXX13 : in std_logic;  
         XXMWX, XFXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX14, 
         MXXXXXXXXXXXXXXXXXXXXX15 : in std_logic);

end XYXX0003;

architecture SYN_USE_DEFA_ARCH_NAME of XYXX0003 is

signal MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, XFXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX3
   , MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX0, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX0, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX1, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX1,
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX2, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX4
   , MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX0, MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX0,
   MXXXXXXXXXXXXXXXXXXXPXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX5, MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWX, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXPXXXXXX10, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX6, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX1, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX3, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXMPXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX1, 
   MXXXXXXXXXXXXXXFXXXXXXXXXX10, MXXXXXXXXXXXXXXFXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX2, 
   MXXXXXXXXXXXXXXFXXXXXXXXXX20, MXXXXXXXXXXXXXXFXXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX3, 
   MXXXXXXXXXXXXXXFXXXXXXXXXX40, MXXXXXXXXXXXXXXFXXXXXXXXXX50, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX4, XFXXXXXXXXXX00, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX5, 
   MXXXXXXXXXXXXXXFXXXXXXXXXX70, XFXXXXXXXXXX20, MXXXXXXXXXXXXXXFXXXXXXXXXXX00,
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXFXXXXXXXXXXX13, MXXXXXXXXXXXXXXFXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXFXXXXXXXXXXX30, MXXXXXXXXXXXXXXFXXXXXXXXXXX40, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXFXXXXXXXXXXX50, MXXXXXXXXXXXXXXFXXXXXXXXXXX60, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX8, 
   MXXXXXXXXXXXXXXFXXXXXXXXXXX70, MXXXXXXXXXXXXXXFXXXXXXXXXXX80, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXFXXXXXXXXXXX90, MXXXXXXXXXXXXXXFXXXXXXXXXXX100, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXFXXXXXXXXXXX110, MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXWXXXXYXX, 
   MXXXXXXXXXXXXXXFXWXXX0, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXVXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXPXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX7, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX8, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX23, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX3, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX0,
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX11, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX12, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX13, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX14, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX16, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX18, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX19, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX20, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX21, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX22, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX23, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX24, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX25, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX26, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX27, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX28, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX29, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX30, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX11, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX12, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXVXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXFXXXXXXXXXXVXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX13, MXXXXXXXXXXXXXXXXXX50, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX14, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXMXMPXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXFXXXHXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX2, MXXXXXXXXXXXXXXXXXXXMXMPXXXX00, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX2, 
   MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX0, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX11
   , MXXXXXXXXXXXXXXXXXXXPXXXX0, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXFXXXHXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXX60, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX, MXXXXXXXXXXXXXXXXXX70, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX0, MXXXXXXXXXXXXXXXXXX80, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX1, MXXXXXXXXXXXXXXXXXX90, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX2, MXXXXXXXXXXXXXXXXXX100, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX
   , MXXXXXXXXXXXXXXXXXX111, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX0, MXXXXXXXXXXXXXXXXXX120, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX1, MXXXXXXXXXXXXXXXXXX130, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX6, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX16, XXMXXXX0_7_port, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXFXXXXXXMXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX17, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX18, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX19, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX7, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX20, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX21, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX22, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX1, 
   MXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX
   , MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX11, MXXXXXXXXXXXXXXXXXXPXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX12, MXXXXXXXXXXXXXXXXXX140, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX23, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX13, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX14, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX24, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX25, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXVXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXX, MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXXXXXFXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX16, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXFXXXXXXXXXXVXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX4, MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX3,
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXX70, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXHXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX32, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX17, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX25, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX6, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXFXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX0, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX1, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX2, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX3, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX4, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX5, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX33, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX0, XXMXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX6, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX34, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX35, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX36, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX37, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX28, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX29, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX31, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX8, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX32, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX33, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX6, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX38, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX39, 
   XXMXXXX0_3_port, XXMXXXX0_6_port, XFXWX0, XXMXXXX0_4_port, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX34, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX3,
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXWXXXXYXX, MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX40,
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX41, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX7, XXMXXXX0_2_port, 
   XXMXXXX0_1_port, MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX35, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX36, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX37, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX9, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX38, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX10, XXMXXXX0_0_port, 
   XXMXXXX0_5_port, MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5, 
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6 : std_logic;

begin
   XFXXXXXXXXXX <= XFXXXXXXXXXX3;
   MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX0;
   MXXXXXXXXXXXXXXXXXXXPXXXXXX <= MXXXXXXXXXXXXXXXXXXXPXXXXXX2;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX <= MXXXXXXXXXXXXXXFXXXXXXXXXXX12;
   MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX1;
   MXXXXXXXXXXXXXXXXXXXPXXXXXX1 <= MXXXXXXXXXXXXXXXXXXXPXXXXXX10;
   MXXXXXXXXXXXXXXFXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXFXXXXXXXXXXXXX0;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX <= 
      MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0;
   MXXXXXXXXXXXXXXFXXXXXXXXXX <= MXXXXXXXXXXXXXXFXXXXXXXXXX10;
   MXXXXXXXXXXXXXXFXXXXXXXXXX1 <= MXXXXXXXXXXXXXXFXXXXXXXXXX11;
   MXXXXXXXXXXXXXXFXXXXXXXXXX2 <= MXXXXXXXXXXXXXXFXXXXXXXXXX20;
   MXXXXXXXXXXXXXXFXXXXXXXXXX3 <= MXXXXXXXXXXXXXXFXXXXXXXXXX30;
   MXXXXXXXXXXXXXXFXXXXXXXXXX4 <= MXXXXXXXXXXXXXXFXXXXXXXXXX40;
   MXXXXXXXXXXXXXXFXXXXXXXXXX5 <= MXXXXXXXXXXXXXXFXXXXXXXXXX50;
   XFXXXXXXXXXX0 <= XFXXXXXXXXXX00;
   MXXXXXXXXXXXXXXFXXXXXXXXXX7 <= MXXXXXXXXXXXXXXFXXXXXXXXXX70;
   XFXXXXXXXXXX2 <= XFXXXXXXXXXX20;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX00;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX1 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX13;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX2 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX20;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX3 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX30;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX4 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX40;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX5 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX50;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX6 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX60;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX7 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX70;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX8 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX80;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX9 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX90;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX10 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX100;
   MXXXXXXXXXXXXXXFXXXXXXXXXXX11 <= MXXXXXXXXXXXXXXFXXXXXXXXXXX110;
   MXXXXXXXXXXXXXXFXWXXX <= MXXXXXXXXXXXXXXFXWXXX0;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX <= 
      MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0;
   MXXXXXXXXXXXXXXXXXXPXXXXXXXX <= MXXXXXXXXXXXXXXXXXXPXXXXXXXX0;
   MXXXXXXXXXXXXXXXXXX5 <= MXXXXXXXXXXXXXXXXXX50;
   MXXXXXXXXXXXXXXXXXXXMXMPXXXX <= MXXXXXXXXXXXXXXXXXXXMXMPXXXX1;
   MXXXXXXXXXXXXXXXXXXXMXMPXXXX0 <= MXXXXXXXXXXXXXXXXXXXMXMPXXXX00;
   MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX <= MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX0;
   MXXXXXXXXXXXXXXXXXXXPXXXX <= MXXXXXXXXXXXXXXXXXXXPXXXX0;
   MXXXXXXXXXXXXXXXXXX6 <= MXXXXXXXXXXXXXXXXXX60;
   MXXXXXXXXXXXXXXXXXX7 <= MXXXXXXXXXXXXXXXXXX70;
   MXXXXXXXXXXXXXXXXXX8 <= MXXXXXXXXXXXXXXXXXX80;
   MXXXXXXXXXXXXXXXXXX9 <= MXXXXXXXXXXXXXXXXXX90;
   MXXXXXXXXXXXXXXXXXX10 <= MXXXXXXXXXXXXXXXXXX100;
   MXXXXXXXXXXXXXXXXXX11 <= MXXXXXXXXXXXXXXXXXX111;
   MXXXXXXXXXXXXXXXXXX12 <= MXXXXXXXXXXXXXXXXXX120;
   MXXXXXXXXXXXXXXXXXX13 <= MXXXXXXXXXXXXXXXXXX130;
   XXMXXXX <= ( XXMXXXX0_7_port, XXMXXXX0_6_port, XXMXXXX0_5_port, 
      XXMXXXX0_4_port, XXMXXXX0_3_port, XXMXXXX0_2_port, XXMXXXX0_1_port, 
      XXMXXXX0_0_port );
   MXXXXXXXXXXXXXXXXXXXXXVXXXXXX <= MXXXXXXXXXXXXXXXXXXXXXVXXXXXX0;
   MXXXXXXXXXXXXXXXXXXPXXXXXX <= MXXXXXXXXXXXXXXXXXXPXXXXXX1;
   MXXXXXXXXXXXXXXXXXX14 <= MXXXXXXXXXXXXXXXXXX140;
   MXXXXXXXXXXXXXXXXXXFXXXXXXX <= MXXXXXXXXXXXXXXXXXXFXXXXXXX0;
   MXXXXXXXXXXXXXXXXXXX7 <= MXXXXXXXXXXXXXXXXXXX70;
   MXXXXXXXXXXXXXXFXXXXXXXXX <= MXXXXXXXXXXXXXXFXXXXXXXXX0;
   XXMXX <= XXMXX0;
   XFXWX <= XFXWX0;
   
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX14, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX,
                           E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           XFXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX0
                           , E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           XFXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX, C 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXXXXX : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX4, C => 
                           MXXXXXXXXXXXXXMXMPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX1 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1, C 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX : MX2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX0 : AX1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX0 : INV port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXX : OR3 port map( A => 
                           MXMXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX3 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX4 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX1 : OR2 port map( A => MXMXXXXXXXXXXXXX, B 
                           => MXMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX2 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX5, A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX6, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX : OA1 port map( A => MXMXXXXXXXXXXXXX0, B
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX1 : OR3A port map( A => 
                           MXMXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX2 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXXXXXX0,
                           C => MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX3 : OR2 port map( A => MXMXXXXXXXXXXXXXXX, B
                           => MXMXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXX1 : OR3B port map( A => 
                           MXMXXXXXXXXXXXXXXXXX0, B => MXMXXXXXXXXXXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXX2 : OR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX4 : OR3 port map( A => MXMXXXXXXXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX4, C => 
                           MXMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXX : OR3 port map( A => MXMXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX3, C => 
                           MXMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX5 : AO13 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXMPXXX, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX5 : OR2 port map( A => MXMXXXXXXXXXXXXX0, B 
                           => MXMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXX2, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, B => 
                           MXMXXXXXXXX, Y => MXXXXXXXXXXXXXXFXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX14, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXXXXX : INV port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX1
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX0, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX1
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX0, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX2 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX1
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX0, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX3 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX2
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX0, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX4 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX2
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX0, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX5 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX3
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX0, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX40);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX6 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX3
                           , E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX50);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX7 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX4
                           , E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           XFXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX8 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX5
                           , E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX9 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX5
                           , E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX70);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX10 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX5
                           , E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           XFXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX11 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX0
                           , E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX7, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX12 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX0
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX13 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX0
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX, Q =>
                           XFXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXX2, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, B => 
                           MXMXXXXXXXX, Y => MXXXXXXXXXXXXXXFXXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX5, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX5, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX6, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX6, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX40);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX7, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX50);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX7, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX60);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX8, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX70);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX8, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX80);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX9, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX90);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX9, Y =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX100);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX10, Y 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX10, Y 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXXX110);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXWXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXWXXXXYXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXFXWXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXVXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXX : OR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX1, B => MXMXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, C => XXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, Y => 
                           XXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXX : INV port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX00, Y => XFXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXWXXXXYXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXWXXXXYXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX4, 
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXXXFX : OR2A port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX10, B => 
                           MXMXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, B => 
                           XFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX60, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX80, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX100, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX110, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX : NOR2B port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX0 : NOR3C port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX1,
                           B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX1, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX1 : OA1A port 
                           map( A => MXMXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX2 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX3, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX3 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX7, 
                           B => MXXXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX4 : NOR3C port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX2,
                           B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX4, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX0, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX5 : NOR3C port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX6, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX6 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX7 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8, 
                           B => XFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX7, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX8 : NOR3C port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX9, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX9 : OA1A port 
                           map( A => MXMXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX10, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX10 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX1, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX11, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX11 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX7, 
                           B => MXXXXXXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX12 : NOR3C port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX12, C 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXMXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX13 : NOR3C port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX14, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX14 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX15 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8, 
                           B => MXXXXXXXXXXXXXXFXXXXXXXXXXX60, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX15, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX16 : OA1A port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXXXXX, C 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX17, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX17 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX18, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX18 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX2, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX19, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX19 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX19);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX20 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8, 
                           B => MXXXXXXXXXXXXXXFXXXXXXXXXXX80, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX20, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX21);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX21 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX22, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX20);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX22 : OA1A port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7
                           , B => MXMXXXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX23, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX22);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX23 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX3, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX23);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX24 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8, 
                           B => MXXXXXXXXXXXXXXFXXXXXXXXXXX100, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX24, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX25);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX25 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX26, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX24);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX26 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX4, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX26);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX27 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8, 
                           B => MXXXXXXXXXXXXXXFXXXXXXXXXXX110, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX27, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX28);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX28 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7
                           , B => MXMXXXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX29, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX27);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX29 : OA1A port 
                           map( A => MXMXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX30, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX29);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXXXX30 : AOI1B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX5, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX30);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX6, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX15, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX0 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXVXXXXXXXXXXXXXXXX : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXVXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXXXXXXX : MX2C port map( 
                           A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXFXXXXXXXXXXVXX
                           , S => MXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXXXX : OA1A port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXX50, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXX : NOR3A port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX1, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXX0 : NOR3B port map( A
                           => MXXXXXXXXXXXXXXXXXXXMXMPXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXFXXXHXXXXXXXXXX, 
                           C => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX2, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXX1 : NOR2B port map( A
                           => MXXXXXXXXXXXXXXXXXXXMXMPXXXX00, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXX2 : OAI1 port map( A 
                           => MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX, C => 
                           MXMXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXXXPXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXFXXX : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXXX50, B => 
                           MXMXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXFXXXHXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXX3 : NOR3B port map( A
                           => MXMXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXX0, C => 
                           MXMXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXX : NOR3C port map( A => 
                           MXMXXXXXXXXXXXXXXX10, B => MXXXXXXXXXXXXXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B =>
                           MXXXXXXXXXXXXXXXXXX60, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX0
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX0 : OA1A port map( A =>
                           XXMXXXXX(3), B => MXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX1, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX1 : OA1A port map( A =>
                           MXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX2 : OA1A port map( A =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B =>
                           MXXXXXXXXXXXXXXXXXX70, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX2, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX3
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX3 : OA1A port map( A =>
                           XXMXXXXX(1), B => MXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX4, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX2
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX4 : OA1A port map( A =>
                           XXXXXXXX, B => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX5 : OA1A port map( A =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B =>
                           MXXXXXXXXXXXXXXXXXX80, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX5, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX6
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX6 : OA1A port map( A =>
                           XXMXXXXX(2), B => MXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX7, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX5
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX7 : OA1A port map( A =>
                           XXXXXXXX0, B => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, C =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX8 : OA1A port map( A =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B =>
                           MXXXXXXXXXXXXXXXXXX90, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX8, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX9
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX9 : OA1A port map( A =>
                           XXMXXXXX(0), B => MXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX10, 
                           Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXXXXXXX10 : OA1A port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXXXXXXX : OA1A port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B
                           => MXXXXXXXXXXXXXXXXXX100, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX, 
                           Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX0)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXXXXXXX0 : AOI1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXXXXXXX1 : OA1A port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B
                           => MXXXXXXXXXXXXXXXXXX111, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX1,
                           Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX2)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXXXXXXX2 : AOI1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX1)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXXXXXXX3 : OA1A port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B
                           => MXXXXXXXXXXXXXXXXXX120, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX3,
                           Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX4)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXXXXXXX4 : AOI1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX3)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXXXXXXX5 : OA1A port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B
                           => MXXXXXXXXXXXXXXXXXX130, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX5,
                           Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX6)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXXXXXXX6 : AOI1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX5)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXXXXXXXXX : AO1D port map( 
                           A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX1 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXFXXXXXXMXXXXXXXXXXXXXXXXX : OR2 port map(
                           A => XXMXXXX0_7_port, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXFXXXXXXMXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX2 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXYXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX3 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXYXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXXXXXX0 : AOI1B port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXX0,
                           C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX5, 
                           Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXXXXXX1 : NOR3B port map( A 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX7, 
                           B => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXXXXXX2 : AOI1 port map( A 
                           => MXXXXXXXXXXXXXXXXXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, B => 
                           XXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, B => 
                           XXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, B => 
                           XXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXXXXXX3 : XA1 port map( A =>
                           MXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXXXXXXX : NOR3B port map( A 
                           => MXXXXXXXXXXXXXXXXXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXX0)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXXXXXVXXXXXXX : OA1 port map(
                           A => MXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXXXXXVXXXXXX : NOR3B port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX
                           , B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX1, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXXXXXVXXXXXX0 : NOR3A port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXPXXXXXXXXLXXXXXLXXVX : OA1 port map(
                           A => MXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXXXXXVXXXXXXX0 : OA1A port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX0, C => 
                           MXXXXXXXXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXPXXXXXXXXLXXXXXLXXVX0 : NOR2B port 
                           map( A => MXXXXXXXXXXXXXXYXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX4 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX11, B => 
                           MXXXXXXXXXXXXXXYXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX11);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX3 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX4 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX3 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX12);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX5 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXXXXXXX : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXX140, B => MXXXXXXXXXXXXXXXXXX15, 
                           C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXXXXXXX1,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXX1)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX, B => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX5 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX : NOR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXX0 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX4 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX14);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX5 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX11, B => XXMXXXX0_7_port, 
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX13);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXXFXX : NOR3B port 
                           map( A => MXXXXXXXXXXXXXXFXWXXX0, B => 
                           XXMXXXX0_7_port, C => XFXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX11, B => XFXXXXXXXXXX00, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXXXXXXXXXXX : NOR3B port map( A =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX24, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX50, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX70, B => XFXXXXXXXXXX00, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXX, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX6 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXXXXXXX : NOR3 port map( 
                           A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXX, Y
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXVXXXXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXVXXXXXXXXXXX, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXVXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, B => 
                           MXMXXXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX4,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, B => 
                           MXMXXXXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX6,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, B => 
                           MXMXXXXXXXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX2,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, B => 
                           MXMXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXXXVXXXXX0,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, B => 
                           MXMXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX0, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, B => 
                           MXMXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX6, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, B => 
                           MXMXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX3, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX, B => 
                           MXMXXXXXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXVXXXXX9, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXX : AO1B port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX28, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX6
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXX0 : AO1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX25, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXX1 : AO1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX21, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX0
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXX2 : AO1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX16, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX5
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXX3 : OR3C port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX1, B =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX13, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX4
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXX4 : AO1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX8, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX2
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXXXXXVXXXXXX1 : OR2 port map(
                           A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX0, B
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX0, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXX0 : OR3C port map( A =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXXXX0, C =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXXFXX0 : NOR3A port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHXXX, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXX1 : NOR3A port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX3, B 
                           => MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX6, B => 
                           XXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXPXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX8, 
                           C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX6, 
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX11);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX1 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX14, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXMXXFXXXXXX : NOR3C port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX25);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXMXXFXXXXXX0 : NOR3B port 
                           map( A => MXXXXXXXXXXXXXXYXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXXFXWXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX2 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX10, Y 
                           => XFXXXXXX(7));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX9, Y =>
                           XFXXXXXX(6));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX8, Y =>
                           XFXXXXXX(5));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX7, Y =>
                           XFXXXXXX(4));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX6, Y =>
                           XFXXXXXX(3));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX6, Y => 
                           XXMXXXXX0(7));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX5, Y => 
                           XXMXXXXX0(6));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX4, Y => 
                           XXMXXXXX0(5));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX3, Y => 
                           XXMXXXXX0(4));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX2, Y => 
                           XXMXXXXX0(3));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX1, Y => 
                           XXMXXXXX0(2));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXX5 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX0, Y => 
                           XXMXXXXX0(0));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX7 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX16);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXMXXX : OR3 port map(
                           A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXX0, 
                           B => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX0, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXFXXXXXXXXXXVXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXVXXXXX5, Y =>
                           XFXXXXXX(2));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXPXXXXXXXXLXXXXXLXXVX1 : AO1B port 
                           map( A => MXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXXXXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXXXXXX,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXPXXXXXXXXLXXXXXLXXVX2 : OR3C port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXX, B => 
                           MXXXXXXXXXXXXXXYXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXX6 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXXVXXXXX, Y => 
                           XXMXXXXX0(1));
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXX5 : AO1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX5, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX1
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXX6 : AO1B port map( A
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXVXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX3
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXX : NOR3A port map( A => 
                           XFXXXXXXXXXX3, B => MXXXXXXXXXXXXXXXXXXFXWXXX2, C =>
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXWXXXXYXXXXXXX0 : NOR3A port map( A => 
                           XXMXXXX0_7_port, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX8, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXWXXXXYXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXX0 : NOR3A port map( A => 
                           XFXXXXXXXXXX00, B => MXXXXXXXXXXXXXXXXXX140, C => 
                           MXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXX140, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXX1, B =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXX2, C =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX24, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX50, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX23);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXFXXX0 : OR3 port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX13, B => 
                           MXMXXXXXXXXXXXXXXX11, C => MXXXXXXXXXXXXXXXXXX50, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXFXXXHXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXX : OR3B port map(
                           A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX0
                           , B => MXXXXXXXXXXXXXXYXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX10, B => 
                           XXXXXXXXXXXXXXXXXX, C => MXXXXXXXXXXXXXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXX70, C => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX12, B => 
                           XXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXXXXX0 : OR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXXXX, C => 
                           MXMXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXX1 : OR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX4, C => 
                           MXMXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX1, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, B => 
                           XXXXXXXX, Y => XFXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX0, Y => 
                           XFXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXX6 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX6 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX2, B => MXXXXXXXXXXXXXXXXXX16, 
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX6 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXX5, Y => MXXXXXXXXXXXXXXXXXXX70
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX8 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXVXXXXXX : OR2 port map( A =>
                           MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXHXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXHXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXX2 : NOR2 port map( A =>
                           MXXXXXXXXXXXXXXXMXMXMXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX9 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX10 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX32, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXFXXXHXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX17);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXXXXXXVXX : OR3A port map( A 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXVXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXFXXXXXXXXXXVXX0, B 
                           => MXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX25);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXFXXXXXXXXXXVXX
                           , B => MXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX23);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXX, B =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX, C => 
                           MXMXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXX : OR3A port map( A => 
                           XXMXXXXX(1), B => MXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7, B => 
                           MXMXXXXXXXXXXXXXXX13, C => MXMXXXXXXXXXXXXXXX14, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXMXXXXXXXX : OR2A port map( 
                           A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXX0 : OR3A port map( A => 
                           XXMXXXXX(3), B => MXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7, B => 
                           MXMXXXXXXXXXXXXXXX15, C => MXMXXXXXXXXXXXXXXX1, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXXXXXXX : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXXX2, A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXX1 : OR3A port map( A => 
                           XXMXXXXX(4), B => MXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXX0 : AO1B port map( A =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7, B => 
                           MXMXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXX2 : OR3A port map( A => 
                           XXMXXXXX(7), B => MXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, C => XXMXXXXX(4), Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, C => XXMXXXXX(5), Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, C => XXMXXXXX(6), Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, C => XXMXXXXX(7), Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXXXX : MX2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXXXX0 : MX2 port map( A => XFXXXXXXXXXXX,
                           S => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, B =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX13, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX30, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX50, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX80, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXXXX5 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX90, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX2 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXMXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXXXXXXX5 : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXXX0 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX1, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX50, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, B => 
                           MXXXXXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXX0 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXXXXXX2, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, B => 
                           MXMXXXXXXXX, Y => MXXXXXXXXXXXXXXFXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXXXXXXX2 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXXXXXXX3 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXVXXXXXX0 : OR2A port map( A 
                           => MXXXXXXXXXXXXXXYXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXX : AOI1 port map( A
                           => MXXXXXXXXXXXXXXXXXXX8, B => MXXXXXXXXXXXXXXXXXXX9
                           , C => MXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXX4 : AOI1 port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX12);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXMXXFXXXXXX1 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXYXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXXXXX : NOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXMXXFXXXXXX2 : NOR3A port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX18, B => 
                           MXXXXXXXXXXXXXXYXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX19);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXMXXFXXXXXX3 : NOR3B port 
                           map( A => MXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX22);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX14 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX0, S => XXMXX0,
                           B => XXMXXXXX(0), Y => MXXXXXXXXXXXXXXXXXX90);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX15 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX1, S => XXMXX0,
                           B => XXMXXXXX(1), Y => MXXXXXXXXXXXXXXXXXX70);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX16 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX2, S => XXMXX0,
                           B => XXMXXXXX(2), Y => MXXXXXXXXXXXXXXXXXX80);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX17 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX3, S => XXMXX0,
                           B => XXMXXXXX(3), Y => MXXXXXXXXXXXXXXXXXX60);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX18 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX4, S => XXMXX0,
                           B => XXMXXXXX(4), Y => MXXXXXXXXXXXXXXXXXX100);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX19 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX5, S => XXMXX0,
                           B => XXMXXXXX(6), Y => MXXXXXXXXXXXXXXXXXX130);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX20 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX6, S => XXMXX0,
                           B => XXMXXXXX(7), Y => MXXXXXXXXXXXXXXXXXX120);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXXFXX1 : AO1 port 
                           map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX34, B => 
                           MXMXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXMXXX0 : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXFXXXXXXXXXXVXX
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXPXXXXXXXXXXXXXXXXXXXXXXXX : NOR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX16);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX33);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXMXXX1 : AO1C port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX21);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXMXXX2 : XAI1A port 
                           map( A => MXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXX4, C => MXXXXXXXXXXXXXXXXXXXXX1,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX20);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXX2 : XA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX17);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX4 : AOI1B port map( A => 
                           MXMXXXXXXXXXXXXXXX16, B => MXMXXXXXXXXXXXXXXX2, C =>
                           MXMXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX36);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX37, B => 
                           MXMXXXXXXXXXXXXXXX17, C => MXMXXXXXXXXXXXXXXX12, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXMXXFXXXXXX4 : NOR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => 
                           MXXXXXXXXXXXXXXYXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXMXXX3 : AO1 port 
                           map( A => MXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX35);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX34, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX1 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX2 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX3 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, B => 
                           XFXXXXXX0(7), C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX4 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX5 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX6 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX7 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX8 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXX0 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, B => 
                           XFXXXXXX0(6), C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX9 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX10 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX11 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX12 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX13 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXX1 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, B => 
                           XFXXXXXX0(4), C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX14 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX15 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXX2 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, B => 
                           XFXXXXXX0(3), C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX16 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX17 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX18 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX19 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX20 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXX3 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, B => 
                           XFXXXXXX0(2), C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX21 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX22 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX23 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX24 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX7, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX25 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX26, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXX4 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, B => 
                           XFXXXXXX0(1), C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX26 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX27 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX28 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX31);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX29 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX32);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX30 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX31, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX33);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXX5 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, B => 
                           XFXXXXXX0(0), C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX90, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX70, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX50, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX30, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX13, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXX5 : MX2 port map( A => XFXXXXXXXXXXX0, S
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXX6 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXXXXXXX4 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXMXXFXXXXXX5 : NOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => 
                           MXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX18);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXWXXPXXXXXXXXXXMXMPXXXXXXXXXXX : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => 
                           MXXXXXXXXXXXXXXYXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXWXXXXYXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXYXX, B => MXXXXXXXXXXXXXXXXXXX12, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX38);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXX0 : XAI1 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX39);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5, B => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7, B => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXPXLXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXX3 : OR3A port map( A => 
                           XXMXXXXX(6), B => MXXXXXXXXXXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXX4 : OR3A port map( A => 
                           XXMXXXXX(5), B => MXXXXXXXXXXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXXXXX : AO1B port map( A 
                           => MXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7, B => 
                           MXMXXXXXXXXXXXXXXX18, C => MXMXXXXXXXXXXXXXXX1, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXX5 : OR3A port map( A => 
                           XXMXXXXX(2), B => MXXXXXXXXXXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXFXXXHX, C => 
                           MXMXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXXXXX2 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXX7, B => 
                           MXMXXXXXXXXXXXXXXX16, C => MXMXXXXXXXXXXXXXXX1, Y =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXXXXXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXXXX1, C 
                           => MXMXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXMXMXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXXXXXXX6 : OR3A port map( A => 
                           XXMXXXXX(0), B => MXXXXXXXXXXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXXFXXXXXXXXXXVXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX4 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX8, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXX1 : XOR2 port map( A => 
                           XXMXXXX0_3_port, B => MXXXXXXXXXXXXXXFXXXXXXXXXX10, 
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXX2 : OR2 port map( A => 
                           XXMXXXX0_6_port, B => MXXXXXXXXXXXXXXXXXXXXXXWXXX, Y
                           => MXXXXXXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXXXXXXXXX : NOR2 port map( A => 
                           XXMXXXX0_3_port, B => MXXXXXXXXXXXXXXFXXXXXXXXXX10, 
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX24);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWXXXXXX0 : NOR2B port map( A => XFXWX0, B
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXWX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXX0 : OR2B port map( A => 
                           XXMXXXX0_6_port, B => XXMXXXX0_4_port, Y => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX5 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXFXXXXXXXXXXXXXXXXX1)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX31 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX32 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX33 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX34 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX34);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9, B => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX6 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX7 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX5 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXHXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXXXXFXWX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXXX4, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXMXMXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX8 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX7 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXXXXFXWX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXXX5, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXWXXXXYXXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXFXXXXXXMXXXXXXXXXXXX, C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXWXXXXYXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXX : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX38, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXYXX, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX40);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXX1 : XO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX41);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXX2 : XA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, C => 
                           MXXXXXXXXXXXXXXYXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX15);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXXXX : XA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX3, C => 
                           MXXXXXXXXXXXXXXYXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXXXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX1, B => MXXXXXXXXXXXXXXXXXXX10
                           , C => MXXXXXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXWXXPXXXXXXXXXXMXMPXXXXXXXXXXX0 : NOR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => 
                           MXXXXXXXXXXXXXXYXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXFXXX1 : OR2A port 
                           map( A => MXMXXXXXXXXXXXXXXX1, B => 
                           MXMXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX13);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX : OR2 port map( A => 
                           MXMXXXXXXXXXXXXXXX1, B => MXMXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXXXX7 : NOR2B port map( A => 
                           MXMXXXXXXXXXXXXX2, B => MXMXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXX5 : NOR2 port map( A 
                           => MXMXXXXXXXXXXXXX0, B => MXMXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXPXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXFXXXXXXXXXX1 : NOR2B port map( A => 
                           XXMXXXX0_2_port, B => XXMXXXX0_1_port, Y => 
                           MXXXXXXXXXXXXXXXXXX140);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXX6 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX31, B => 
                           XFXXXXXX0(5), C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX35 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX34, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX35);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX36 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX9, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX9, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX38, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX37);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX37 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX36);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXVXXXXX38 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX0, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXX38);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXXXX21 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX7, S => XXMXX0,
                           B => XXMXXXXX(5), Y => MXXXXXXXXXXXXXXXXXX111);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXMXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11, B => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXMXXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXXXMXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX9 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXXX6, B => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXLXXMXXX10);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXPXXXXXXXXXXMXMPXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXX3 : OR3B port map( A =>
                           MXMXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXX4, C => 
                           MXMXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXMXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXXXXXXX : NOR2B port 
                           map( A => MXMXXXXXXXXXXXXX5, B => MXMXXXXXXXXXXXXX4,
                           Y => MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXXXXX : NOR3B port map(
                           A => MXMXXXXXXXXXXXXX2, B => MXMXXXXXXXXXXXXX, C => 
                           MXMXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXXFXX2 : OR3B port 
                           map( A => MXMXXXXXXXXXXXXX6, B => MXMXXXXXXXXXXXXX5,
                           C => MXMXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX34);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXFXXX2 : OR3C port 
                           map( A => MXMXXXXXXXXXXXXX6, B => MXMXXXXXXXXXXXXX5,
                           C => MXMXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX37);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXFXXX3 : OR3B port 
                           map( A => MXMXXXXXXXXXXXXX3, B => MXMXXXXXXXXXXXXX0,
                           C => MXMXXXXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXXXX50);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXXXXXXX0 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXYXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXFXXX4 : NOR3A port 
                           map( A => MXMXXXXXXXXXXXXX3, B => MXMXXXXXXXXXXXXX, 
                           C => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX14);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXPXXXXXXXXXXXXFXXX5 : AOI1 port 
                           map( A => MXMXXXXXXXXXXXXX6, B => MXMXXXXXXXXXXXXX5,
                           C => MXXXXXXXXXXXXXXXXXX50, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX32);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXXXXX0 : OR2A port map(
                           A => MXMXXXXXXXXXXXXX, B => MXMXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX00);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXPXXXXXXXXXXMXMPXXXXXX6 : OA1B port map( C 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX3, A => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXPXXXXXXXXXXXXXXVXXX : AO1C port map( A 
                           => MXXXXXXXXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX, C =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXVXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXX3 : XAI1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, C => 
                           MXXXXXXXXXXXXXXYXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX11 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXX9, C => XXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX12 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXXXXXX13 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX9, B => MXXXXXXXXXXXXXXXXXX25,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX15);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXX26, B => MXXXXXXXXXXXXXXXXXX21, Y
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXPXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX7, CLK =>
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXLXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXHXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXMXMPXXXXXX6, CLK =>
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXPXHXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXVXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLXXVXXX, CLK =>
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXWXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXWXXXXYXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => XFXWX0
                           );
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMWXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXWXXXXYXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => XXMWX)
                           ;
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXXXVXXXX, E => 
                           MXXXXXXXXXXXXXMXMPXXXXX, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Q => XXMXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXFXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXMXMPXXXXXXXX, E => 
                           MXXXXXXXXXXXXXMXMPXXXXX, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, Q => XFXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXX : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX0, CLK => XLXXPX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXX0 : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX1, CLK => XLXXPX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXX1 : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX2, CLK => XLXXPX, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX3, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX4, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXXX1, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX5, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX6, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXPXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXX2 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q =>
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXX3 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXX4 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXX5 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX0, E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXXXX6 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXYXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXXXVXXXXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX1
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXX0, Q 
                           => XXMXXXX0_0_port);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXX0 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX2
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX15, Q =>
                           XXMXXXX0_1_port);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX3
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX15, Q =>
                           XXMXXXX0_2_port);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXX2 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX4
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX15, Q =>
                           XXMXXXX0_3_port);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXX3 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX5
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX15, Q =>
                           XXMXXXX0_4_port);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXX4 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX0
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX15, Q =>
                           XXMXXXX0_5_port);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXX5 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX,
                           E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, CLK
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX15, Q => 
                           XXMXXXX0_6_port);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXFXXXXXXXX6 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXMXXFXXXXXXXXXXXXYXXXXX6
                           , E => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX22, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXXXXXX, Q 
                           => XXMXXXX0_7_port);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX2 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX, C 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX3 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, C 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX4 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, C 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, Y 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX6 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX7 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3, B 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXMPXXX,
                           Y => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX8 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX9 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX10 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6, B 
                           => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX11 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX12 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX13 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX14 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX15 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX16 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX17 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX18 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX19 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX20 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXXX21 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2);
   MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXXX3 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXPXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXWXXXXXXXXXXXXXXMPXXX);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity XYXX0002 is

   port( MXXXXXXXXXXXXXXXXXXXFXWXXX, MXXXXXXXXXXXXXXXXXXFXWXXX : out std_logic;
         MXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, XLXXPX, MXXXXXXXXXXXXXXXXXXXXXXXX : 
         in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX : out std_logic;  ramaddr : in 
         std_logic_vector (4 downto 2);  XFXXXXXXXXXX, XFXXXXXXXXXXXX : in 
         std_logic;  MXXXXXXXXXXXXXXXXXXFXWXXX0 : out std_logic;  
         MXXXXXXXXXXXXXXYXX, MXXXXXXXXXXXXXMXMPXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXX
         , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX, MXXXXXXXXXXXXXMXMPXXXXXX : 
         in std_logic;  MXMPXXXXWXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXYXXXXXX, 
         MXXXXXXXXXXXXXMXMPXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX0 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXFXWXXXXX : out 
         std_logic;  MXXXXXXXXXXXXXXXXXXXX : in std_logic;  MXMPXXX : out 
         std_logic;  XFXXXXXXXXXX0, XFXXXXXXXXXX1 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXFXWXXXXX : out std_logic;  XXXXXPXXX : in std_logic
         ;  MXXXXXXXXXXXXXXXMXMXXXLXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXYXXXX, MXXXXXXXXXXXXXXXXXXXXXXXVXX, 
         MXXXXXXXXXXXXXXXXXFXXXHX, MXXXXXXXXXXXXXXXXXXLLXX, 
         MXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX0, 
         MXXXXXXXXXXXXXPXLXXXXXX1 : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX1 : 
         in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX2 : out std_logic;  XXXXXXXX : 
         in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX3 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXX2 : in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX4 : 
         out std_logic;  XXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXX3 : in std_logic;  
         MXXXXXXXXXXXXXPXHXXXXXX, MXXXXXXXXXXXXXPXHXXXXXX0 : out std_logic;  
         MXMXXXX : out std_logic_vector (15 downto 0);  XXXXXXXX1, XXXXXXXX2, 
         MXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXXXVXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXXXVXXXXXX2, MXXXXXXXXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXXXVXXXXXX3, MXXXXXXXXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXPXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXX4, MXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXHXXX, MXXXXXXXXXXXXXXXXXXXHXXX0, 
         MXXXXXXXXXXXXXXXXXXXHXXX1, MXXXXXXXXXXXXXXXXXXXXX4, 
         MXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX6, XXXXXXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXX7, MXMXXXX0, MXXXXXXXXXXXXXXXXXXX8, 
         MXXXXXXXXXXXXXXXXVXLXX, MXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXX10,
         MXXXXXXXXXXXXXXYXXXX0, MXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXX12,
         MXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXXXXXX2 : in std_logic;  
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2, 
         MXXXXXXXXXXXXXXXXXXFXXXXXXX, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9, 
         MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11
         , MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12 : out std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXWXXX, 
         MXXXXXXXXXXXXXXFXWXXX : in std_logic;  XXMXXXXX : in std_logic_vector 
         (7 downto 0);  MXXXXXXXXXXXXXXFXXXXXMXXXXX : out std_logic;  
         MXMXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXX0 : in std_logic;  
         MXXXXXXXXXXXXXPXHXXXXXX1, MXXXXXXXXXXXXXPXHXXXXXX2, 
         MXXXXXXXXXXXXXPXHXXXXXX3, MXXXXXXXXXXXXXPXHXXXXXX4, 
         MXXXXXXXXXXXXXPXLXXXXXX5 : out std_logic;  MXXXXXXXXXXXXXXXXXXFXWXXX1,
         MXMXXXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXXXX3 : in 
         std_logic;  MXXXXXXXXXXXXXPXHXXXXXX5, MXXXXXXXXXXXXXPXHXXXXXX6, 
         MXXXXXXXXXXXXXPXLXXXXXX6 : out std_logic;  MXXXXXXXXXXXXXXYXX0, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXX0, MXXXXXXXXXXXXXMXMPXXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXJXMP, MXXXXXXXXXXXXXXXXXXX15 :
         in std_logic;  MXXXXXXXXXXXXXXXXXMXVXWXXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXMXMPXXXXXXX2, 
         MXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXXXXXFXWXXX2 : 
         out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXWXXX0, MXMXXXXXXXXXXXXXXX4, 
         MXMXXXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXFXXXHX : 
         in std_logic;  MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX : out 
         std_logic;  MXXXXXXXXXXXXXXYXXXX1, MXXXXXXXXXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXLL : in std_logic;  MXMXXXXX : in std_logic_vector 
         (7 downto 0);  MXMXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXXXPXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, XFXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX5, MXXXXXXXXXXXXXXFXXXXXXXXX, 
         MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX9, MXMXXXXXXXXXXXXXXX10, 
         MXMXXXXXXXXXXXXXXX11, MXMXXXXXXXXXXXXXXX12, MXMXXXXXXXXXXXXXXX13, 
         MXMXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXYFLXX, 
         MXXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXYXX1 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXPXXLXX : out std_logic;  MXXXXXXXXXXXXXXXXXXX20, 
         MXXXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXX4, XXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXXXX15, MXMXXXXXXXXXXXXXXX16, 
         MXMXXXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX5 : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXFXWXXX0 : out std_logic;  XFXWX, 
         MXXXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXMXMPXXXX : out
         std_logic;  MXXXXXXXXXXXXXXXXXXX21, XXMXXXXXXX, 
         MXXXXXXXXXXXXXMXMPXXXXX, XXXXXXXX3, MXXXXXXXXXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXXXXFXXXHXXX, MXXXXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXX6 : in std_logic;  
         MXXXXXXXXXXXXXXXMXMXMXXXX, MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, 
         MXMWXXXXXX, MXXXXXXXXXXXXXMXMXXXX, MXMXX : out std_logic;  XFXXXXXX : 
         in std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXXXXXXXXX7, 
         MXMXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXX3, 
         MXMXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXX6, 
         MXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXX9, 
         MXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXX11, 
         MXXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXXX13, 
         MXXXXXXXXXXXXXXXXXXXXX14 : in std_logic);

end XYXX0002;

architecture SYN_USE_DEFA_ARCH_NAME of XYXX0002 is

signal MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX0, MXXXXXXXXXXXXXXXXXXXFXWXXX1, 
   MXXXXXXXXXXXXXXXXXXFXWXXX3, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMMX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, MXXXXXXXXXXXXXPXLXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX4, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX9, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX6, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0, 
   MXXXXXXXXXXXXXXXXXXFXWXXX00, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXL, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, MXMPXXXXWXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX3, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX6,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, MXXXXXXXXXXXXXXXXXXFXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX10, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX
   , MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWX, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXX, MXXXXXXXXXXXXXPXLXXXXXX00, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX, MXXXXXXXXXXXXXPXLXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX10, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX2, MXXXXXXXXXXXXXPXLXXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX1, MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX3
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX3, MXXXXXXXXXXXXXPXLXXXXXX30, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX18, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX4, MXXXXXXXXXXXXXPXLXXXXXX40, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX22, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX3, MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX5
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX23, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX24, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX5, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX25, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX26, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX27, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX28, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX, MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX1
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX6, MXXXXXXXXXXXXXPXHXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX3, MXXXXXXXXXXXXXPXHXXXXXX00, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX8, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX29, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX30, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX31, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX32, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX33, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX34, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX35, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX36, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXX,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX37, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX38, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX39, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX40, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX19, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX22
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX20, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX21, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX22, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX23, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX24, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX25, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX28, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX26, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX27, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX28, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX29, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX30, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX31, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX32, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX33, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX34, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX31, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX32, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX2, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX35
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX33, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX4, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX36
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX34, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX6, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX37
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX35, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX8, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX38
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX36, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX39, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX4, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX37,
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX40, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX38, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX41, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX29, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX42, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX43, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX44, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX45, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX46, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX47, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX48, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX4, 
   MXMXXXX1_0_port, MXMXXXX1_1_port, MXMXXXX1_2_port, MXMXXXX1_3_port, 
   MXMXXXX1_4_port, MXMXXXX1_5_port, MXMXXXX1_6_port, MXMXXXX1_7_port, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX2, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX3, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX4, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX5, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX6, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX6, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX49, MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX0
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX2, MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX3, MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX4, MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX5, MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX1
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXFFXXLXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL0
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX0,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX2, MXXXXXXXXXXXXXXXMXMXXXLXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXWXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXMMX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX0, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX13, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX5, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16,
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX6, 
   MXXXXXXXXXXXXXXXXXXFXXXXXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX2, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX3, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX4, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX5, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX2, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX4, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX2, MXMXXXX1_11_port, 
   MXMXXXX1_10_port, MXMXXXX1_9_port, MXMXXXX1_8_port, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX39, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX28, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX40, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX29, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX41, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX42, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX31, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX43, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX31, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX20
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX32, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX21, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX33
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX22, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX34, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX23
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX35, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX24, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX36
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX25, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX37, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX26
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX38, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX27, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX39
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX28, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX40, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX29
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX41, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX42, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX43, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX44, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX45, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX46, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX32, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX44, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX33, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX45
   , MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX34, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX46, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX35, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX47, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX36, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX48, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX37, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX49, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX38, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX50, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX39, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX51, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX40, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX52, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX41, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX53, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX14, MXXXXXXXXXXXXXPXHXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2, MXXXXXXXXXXXXXPXHXXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX16, MXXXXXXXXXXXXXPXHXXXXXX30, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX3, MXXXXXXXXXXXXXPXHXXXXXX40, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX39, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX40, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX41, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX42, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX43, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX44, MXXXXXXXXXXXXXPXLXXXXXX50, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX45, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX6, MXXXXXXXXXXXXXPXHXXXXXX50, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX7, MXXXXXXXXXXXXXPXHXXXXXX60, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX46, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX47, MXXXXXXXXXXXXXPXLXXXXXX60, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX48, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX49, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX50, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX51, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX52, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX53, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX54, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX55, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX2, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL4, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXXLX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX2
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX50, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX51, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX3, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, MXXXXXXXXXXXXXXXXXXFXWXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX42, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX54, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXHXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX1,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX6, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX7, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX8, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX9, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX10, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX11, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX12, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX2
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX21
   , MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXMXMXXXLXMXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXX1, MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX41, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX42, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX43, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX44, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, MXMXXXX1_12_port, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, MXMXXXX1_13_port, MXMXXXX1_14_port, 
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12, MXMXXXX1_15_port, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX22, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXXXX
   , MXXXXXXXXXXXXXXXMXMXXXLXMXVXXXXFF, MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX3, MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX5, MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX6, 
   MXXXXXXXXXXXXXXXXXXXFXWXXX00, MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX2, 
   MXXXXXXXXXXXXXXXXXXMXMPXXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX3,
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX12, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX53, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX54, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX55, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX56, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX57, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX58, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX59, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX60, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX61, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX62, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX63, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX64, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX65, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX66, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX67, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX8, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX10, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX12, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX14, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX16, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX18, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX20, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX0, MXXXXXXXXXXXXXXXMXMXXXLXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXX1, MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXX2, MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXXXX3, MXXXXXXXXXXXXXXXMXMXXXLXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX19, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX7, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX8, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX9, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX0, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX10, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX1, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX11, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX2, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX12, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX13, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX14, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX3, 
   MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX4 : std_logic;

begin
   MXXXXXXXXXXXXXXXXXXXFXWXXX <= MXXXXXXXXXXXXXXXXXXXFXWXXX1;
   MXXXXXXXXXXXXXXXXXXFXWXXX <= MXXXXXXXXXXXXXXXXXXFXWXXX3;
   MXXXXXXXXXXXXXPXLXXXXXX <= MXXXXXXXXXXXXXPXLXXXXXX7;
   MXXXXXXXXXXXXXXXXXXFXWXXX0 <= MXXXXXXXXXXXXXXXXXXFXWXXX00;
   MXMPXXXXWXXX <= MXMPXXXXWXXX0;
   MXXXXXXXXXXXXXXXXXXFXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXFXXXXXXXXX0;
   MXXXXXXXXXXXXXXXXXXXFXWXXXXX <= MXXXXXXXXXXXXXXXXXXXFXWXXXXX0;
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX <= MXXXXXXXXXXXXXXXMXMXXXLXXXXXX10;
   MXXXXXXXXXXXXXPXLXXXXXX0 <= MXXXXXXXXXXXXXPXLXXXXXX00;
   MXXXXXXXXXXXXXPXLXXXXXX1 <= MXXXXXXXXXXXXXPXLXXXXXX10;
   MXXXXXXXXXXXXXPXLXXXXXX2 <= MXXXXXXXXXXXXXPXLXXXXXX20;
   MXXXXXXXXXXXXXPXLXXXXXX3 <= MXXXXXXXXXXXXXPXLXXXXXX30;
   MXXXXXXXXXXXXXPXLXXXXXX4 <= MXXXXXXXXXXXXXPXLXXXXXX40;
   MXXXXXXXXXXXXXPXHXXXXXX <= MXXXXXXXXXXXXXPXHXXXXXX7;
   MXXXXXXXXXXXXXPXHXXXXXX0 <= MXXXXXXXXXXXXXPXHXXXXXX00;
   MXMXXXX <= ( MXMXXXX1_15_port, MXMXXXX1_14_port, MXMXXXX1_13_port, 
      MXMXXXX1_12_port, MXMXXXX1_11_port, MXMXXXX1_10_port, MXMXXXX1_9_port, 
      MXMXXXX1_8_port, MXMXXXX1_7_port, MXMXXXX1_6_port, MXMXXXX1_5_port, 
      MXMXXXX1_4_port, MXMXXXX1_3_port, MXMXXXX1_2_port, MXMXXXX1_1_port, 
      MXMXXXX1_0_port );
   MXXXXXXXXXXXXXXXXXXFXXXXXXX <= MXXXXXXXXXXXXXXXXXXFXXXXXXX0;
   MXXXXXXXXXXXXXPXHXXXXXX1 <= MXXXXXXXXXXXXXPXHXXXXXX10;
   MXXXXXXXXXXXXXPXHXXXXXX2 <= MXXXXXXXXXXXXXPXHXXXXXX20;
   MXXXXXXXXXXXXXPXHXXXXXX3 <= MXXXXXXXXXXXXXPXHXXXXXX30;
   MXXXXXXXXXXXXXPXHXXXXXX4 <= MXXXXXXXXXXXXXPXHXXXXXX40;
   MXXXXXXXXXXXXXPXLXXXXXX5 <= MXXXXXXXXXXXXXPXLXXXXXX50;
   MXXXXXXXXXXXXXPXHXXXXXX5 <= MXXXXXXXXXXXXXPXHXXXXXX50;
   MXXXXXXXXXXXXXPXHXXXXXX6 <= MXXXXXXXXXXXXXPXHXXXXXX60;
   MXXXXXXXXXXXXXPXLXXXXXX6 <= MXXXXXXXXXXXXXPXLXXXXXX60;
   MXXXXXXXXXXXXXXXXXXFXWXXX2 <= MXXXXXXXXXXXXXXXXXXFXWXXX20;
   MXXXXXXXXXXXXXXXXXXXFXWXXX0 <= MXXXXXXXXXXXXXXXXXXXFXWXXX00;
   MXXXXXXXXXXXXXXXXXXMXMPXXXX <= MXXXXXXXXXXXXXXXXXXMXMPXXXX0;
   
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXFFXXXXXXXXXFXWXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMMX, B => 
                           MXXXXXXXXXXXXXXXXXXX, C => MXXXXXXXXXXXXXXXXXXXXX, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMMX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX3 : OR2 port map( A => ramaddr(3), B => 
                           ramaddr(4), Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX1 : NOR3 port map( A => XFXXXXXXXXXX, B => 
                           XFXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX00);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX2 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX3 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX4 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMMX, B => 
                           MXXXXXXXXXXXXXXXXXXX, C => MXXXXXXXXXXXXXXXXXXXXX, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXL);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX : AX1D port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX,
                           B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0
                           );
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX1 : MAJ3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX)
                           ;
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX2 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX
                           , B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX4 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0
                           , B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX0, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX1
                           );
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX1
                           , B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX
                           );
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX5 : AO1B port map( A => MXXXXXXXXXXXXXXYXX, B 
                           => MXXXXXXXXXXXXXMXMPXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMMX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX6 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXX, Y => MXMPXXXXWXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX7 : OR2 port map( A => XFXXXXXXXXXXXX, B => 
                           XFXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXXXXFXWXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX0, B => MXXXXXXXXXXXXXXXXXXXXXX0
                           , C => MXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX, B => 
                           MXXXXXXXXXXXXXXYXXXXXX, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX, B => 
                           MXXXXXXXXXXXXXXYXXXXXX, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXXXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXXXXX1 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXXXXXXX0 : OA1B port map( C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMMX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXXXXX : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX5, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX5 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX6 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX7 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX8 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX9 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX4, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX10 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX11 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX5, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX12 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX7, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX5, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX0, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX5 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX6 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX3, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX7 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX8 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX6, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX9 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX4, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX10 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX10, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX11 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX7, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX12 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMPXXXXX : INV port map( A => MXMPXXXXWXXX0, Y => 
                           MXMPXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX : NOR2 port map( A => XFXXXXXXXXXX0, B 
                           => XFXXXXXXXXXX1, Y => MXXXXXXXXXXXXXXXXXXFXWXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXXXXX : NOR2A port map( A => XXXXXPXXX,
                           B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXXXXXXX : NAND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWXXXXXX0 : NAND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, B => 
                           MXXXXXXXXXXXXXXXXXXLLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXX : NAND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXX0 : NAND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWX, B => 
                           MXXXXXXXXXXXXXXXXXXLLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX4 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX6, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX6 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX11 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX12 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX13 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX14 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX15 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX16 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, B => 
                           XXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX17 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX18 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX19 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX20 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX21 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX22 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX23 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX5, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX24);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX24 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, B => 
                           XXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX23);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX25 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX26);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX26 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX27);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX27 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX6, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX25);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX28 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX28);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX5, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX6, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX29 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX29);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX30 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX30);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX31 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX31);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX32 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX32);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX33 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX33);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX34 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX34);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX35 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX35);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX36 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX36);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX37 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX37);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXX38 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX38);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXXX3 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX39, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXXXXXXX4 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX19, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX7 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX25, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX9 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX26, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX11 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX27, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX12 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX13 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX28, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX14 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX15 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX16 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX17 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXX18 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX28, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX29, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX32, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX7 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX33, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX9 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX34, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX31, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX32, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX34, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX7 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX35, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX9 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX36, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX39, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX11 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX12 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX13 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX14 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX41, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX15 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX29, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX16 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX42, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX17 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXX18 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX44, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX45, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX46, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX7 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX25, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX47, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX9 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX26, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX48, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXXX : NOR2A port map( A => 
                           MXMXXXX1_0_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXXX0 : NOR2A port map( A => 
                           MXMXXXX1_1_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXXX1 : NOR2A port map( A => 
                           MXMXXXX1_2_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXXX2 : NOR2A port map( A => 
                           MXMXXXX1_3_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXXX3 : NOR2A port map( A => 
                           MXMXXXX1_4_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXXX4 : NOR2A port map( A => 
                           MXMXXXX1_5_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXXX5 : NOR2A port map( A => 
                           MXMXXXX1_6_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXXX6 : NOR2A port map( A => 
                           MXMXXXX1_7_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXXXXXXX0 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, B => 
                           XXXXXXXX1, C => MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX1, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXXXXXXX1 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXLXX, B => 
                           XXXXXXXX2, C => MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX2, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXXXXXXX2 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXL, B => 
                           MXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXXXXXXX3 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXL, B => XXXXXXXX,
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXXXXXXX4 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXL, B => 
                           MXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXXXXXXX5 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXL, B => XXXXXXXX0
                           , C => MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXXXXXXX6 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXL, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXLLXX, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX49, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX1 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXLLXX, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX4 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXLLXX, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX6 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX7 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX8 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXLLXX, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX1, B => MXXXXXXXXXXXXXXXXXXXX, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX10 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXXXX11 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXLLXX, B => 
                           MXXXXXXXXXXXXXXXXVXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX3, B => MXXXXXXXXXXXXXXXXXXXXX, 
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX0, B => 
                           MXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXXXXXXX1 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => MXXXXXXXXXXXXXXXXXFXXXHX
                           , C => MXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXXXXXXXXX : OA1A port map( A =>
                           MXXXXXXXXXXXXXXXXXXXHXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXMXXX, Y =>
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXXXXXXXXX0 : OA1A port map( A 
                           => MXXXXXXXXXXXXXXXXXXXHXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXMXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXVXXXXXXXXXX : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX3, S => 
                           MXXXXXXXXXXXXXXXXXXXHXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXFFXXLXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXX6, A => XXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXWXXXXXXXXXX : NOR2 port map( A => MXMXXXX0,
                           B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXWXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX8, B => MXXXXXXXXXXXXXXXXVXLXX, 
                           C => MXXXXXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXFFXXLXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX8, B => MXXXXXXXXXXXXXXXXXXX10, 
                           C => MXXXXXXXXXXXXXXYXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXFFXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXMXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXXXXXXX2 : NOR2B port map( A => MXMXXXX0, 
                           B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXMMX, B => 
                           MXXXXXXXXXXXXXXYXXXX0, C => MXXXXXXXXXXXXXXXXXXXX, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL, B => 
                           MXXXXXXXXXXXXXXYXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMX0, B => 
                           MXXXXXXXXXXXXXXYXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXVXLXX, B => MXXXXXXXXXXXXXXXXXXX12,
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXXXXXXX2 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX, B => MXXXXXXXXXXXXXXXXXXXXXXX2
                           , Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXMMX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX13, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX, B => XFXXXXXXXXXX1, 
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX14, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX0, B => XFXXXXXXXXXX1,
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX9, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX1, B => XFXXXXXXXXXX1,
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX3, B => 
                           XFXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX5 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX10, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX18, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX2, B => XFXXXXXXXXXX1,
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX19, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX3, B => XFXXXXXXXXXX1,
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX20, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX4, B => XFXXXXXXXXXX1,
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX11 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX12 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX21, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXXXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX5, B => XFXXXXXXXXXX1,
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXFFXXXXXXXXXFXWXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, B => XFXXXXXXXXXX1, C 
                           => MXXXXXXXXXXXXXXXXXXXXXXWXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXFXWXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXWXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXX0, C => XXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX1, B => XXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX2, B => XXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX3, B => XXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXX : OR3B port map( A => 
                           MXMXXXX1_11_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXX0 : OR3B port map( A => 
                           MXMXXXX1_10_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXX1 : OR3B port map( A => 
                           MXMXXXX1_9_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXX2 : OR3B port map( A => 
                           MXMXXXX1_8_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0, B => 
                           XXMXXXXX(7), C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0, B => 
                           XXMXXXXX(6), C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0, B => 
                           XXMXXXXX(5), C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0, B => 
                           XXMXXXXX(4), C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0, B => 
                           XXMXXXXX(3), C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXX4 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0, B => 
                           XXMXXXXX(2), C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXX5 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0, B => 
                           XXMXXXXX(1), C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXX6 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0, B => 
                           XXMXXXXX(0), C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX0, B => 
                           XXXXXXXXXXXXXXXX, C => MXXXXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX12, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXFXXXXXMXXXXVXXXXX17, Y => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, B => 
                           MXMXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, B => 
                           MXMXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX39);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX28, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX40);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXX1 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX29, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX41);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXX2 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX42);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXX3 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX43);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX32, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX1 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX33, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX2 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX34, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX23);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX3 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX24);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX25);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX5 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX26);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX6 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX27);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX7 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX39, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX28);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXX8 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX29);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX41);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX42);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXX1 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX43);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXX2 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX44);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXX3 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX45);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX46);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX32, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX44);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX33, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX45);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX1 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX34, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX46);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX2 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX47);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX3 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX48);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX49);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX5 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX50);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX6 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX39, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX51);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX7 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX52);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXX8 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX41, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX53);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX27, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX39);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX24, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX40);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX20, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX41);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX16, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX5, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX42);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX6, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX43);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX4 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX44);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX5 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX50, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX45);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX00, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, B => 
                           MXMXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, B => 
                           MXMXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXXXXX0 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, B => 
                           MXMXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX50, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX60, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX6 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX38, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX46);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX7 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX47);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX8 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX60, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX48);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX9 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX49);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX10 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX30, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX50);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX11 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX33, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX51);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX12 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX52);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX13 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX00, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX31, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX53);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX14 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX54);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXX15 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX50, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX55);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXYXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX13 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => MXXXXXXXXXXXXXXXJXMP, C
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXWXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL0, B => MXMXXXX0, C
                           => MXXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXMXVXWXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL4, C => 
                           MXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL1, B => 
                           MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXFFXXXXXXXXXFXWX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXXLX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXHXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXHXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXX0 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL, C => 
                           MXXXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXX2 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => MXXXXXXXXXXXXXXXXXXXX0,
                           C => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXX0 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX14 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX0, B => MXXXXXXXXXXXXXXXXXXXX0, 
                           C => MXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXVXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXVXXXXX, C 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXMXXX, 
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX50, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXXXX0, 
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX51, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXXXX, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXX3 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMMX, C => 
                           MXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX00, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX00, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX00, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, B => 
                           MXMXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXXX2 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX42, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXVXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX54);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, B => 
                           MXMXXXXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0, B => 
                           MXMXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXHXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX, C => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXYXXXX1, B => MXXXXXXXXXXXXXXXXXXX6, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX6, B => MXXXXXXXXXXXXXXXXXXXX1, 
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXYXXXX1, B => MXXXXXXXXXXXXXXXXXXX17, 
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWXXXXXX1 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXLLXX, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFLWXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMMX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX0 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX1 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX2 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX3 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX4 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX5 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX6 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX7 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX8 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX9 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX10 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX11 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX12 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX13 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX14 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX15 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXVXXXXX6, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX16 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX7, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX0 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX1 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX2 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX3 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX4 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX5 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX0, C => 
                           MXXXXXXXXXXXXXXYXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXLLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX0 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXLLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXLL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX0 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXLL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX1 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXLL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX2 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXLL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX3 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX10, C =>
                           MXXXXXXXXXXXXXXXXXXLL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX4 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXVXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXXLL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXXXXX : NOR2A port map( A => MXMXXXXX(1),
                           B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXXXXX0 : NOR2A port map( A => MXMXXXXX(2)
                           , B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXXXXX1 : NOR2A port map( A => MXMXXXXX(3)
                           , B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXXXXX2 : NOR2A port map( A => MXMXXXXX(4)
                           , B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXXXXX3 : NOR2A port map( A => MXMXXXXX(5)
                           , B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXXXXX4 : NOR2A port map( A => MXMXXXXX(6)
                           , B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX : NOR2A port map( A => MXMXXXXX(7), B =>
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX5 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXX7 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX42, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX43, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX44, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXXXXXXX : OR2B port map( A => MXMXXXXX(1)
                           , B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, Y =>
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXXXXXXX0 : OR2B port map( A => 
                           MXMXXXXX(2), B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX60, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXX5 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXX5 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXHXXXXXX60, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXX1 : OR2B port map( A => 
                           MXMXXXX1_12_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXPXHXXXXXX50, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXPXXMXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXX2 : OR2B port map( A => 
                           MXMXXXX1_13_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXX3 : OR2B port map( A => 
                           MXMXXXX1_14_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXXXXXXX4 : OR2B port map( A => 
                           MXMXXXX1_15_port, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXMXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXMXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX4 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXLXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX5 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX6 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX7 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX42, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX43, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX44, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXXX4 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX40, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX5 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX7 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX8 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX5 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX7 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX8 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXXXXXXX : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX : OR2B port map( A => 
                           XXMXXXXX(3), B => MXXXXXXXXXXXXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX0 : OR2B port map( A => 
                           XXMXXXXX(7), B => MXXXXXXXXXXXXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXXXMXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, B => 
                           XXMXXXXX(1), Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX1 : OR2B port map( A => 
                           XXMXXXXX(2), B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX2 : OR2B port map( A => 
                           XXMXXXXX(6), B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX3 : OR2B port map( A => 
                           XXMXXXXX(7), B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX9 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX9 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX10 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXX10 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX11 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX4 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXX12 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX5 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX5 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX6 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX7 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX7 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX8 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX8 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX9 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX : MX2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX40);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX0 : MX2C port map( A => XFXXXXXXXXXXX, S 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX39);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX38);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX37);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX3 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX36);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX4 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX35);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX5 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX34);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX6 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX33);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX7 : MX2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX32);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX8 : MX2C port map( A => XFXXXXXXXXXXX, S 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX31);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX31);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX0 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX3 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX4 : MX2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX41);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX5 : MX2C port map( A => XFXXXXXXXXXXX, S 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX40);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX6 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX39);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX7 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX38);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX8 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX37);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX9 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX36);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX10 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX35);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX11 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX34);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX12 : MX2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX33);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX13 : MX2C port map( A => XFXXXXXXXXXXX, S
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX32);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX0 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX3 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX4 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX14 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19, B => 
                           MXMXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX15 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19, B => 
                           MXMXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX5 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX19, B => 
                           MXMXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX6 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX7 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX8 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX9 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX10 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXMXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX3 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX4 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX5 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX6 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXX7 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX41);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX0 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX42);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX43);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX44);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX3 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX39);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXX4 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX40);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX : MX2C port map( A => MXMXXXXXXXXXXXXXXX8,
                           S => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX31);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX0 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX32);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX1 : MX2C port map( A => MXMXXXXXXXXXXXXXXX9
                           , S => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX33);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX2 : MX2C port map( A => MXMXXXXXXXXXXXXXXX7
                           , S => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX34);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX3 : MX2C port map( A => MXMXXXXXXXXXXXXXXX4
                           , S => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX35);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX4 : MX2C port map( A => MXMXXXXXXXXXXXXXXX6
                           , S => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX36);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX5 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX37);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX6 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX38);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX9 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX10 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX11 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX12 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX13 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX14 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX15 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX16 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX16 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX17 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX18 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX13, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX19 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX20 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXMXMXXXLXMX : MX2 port map( A => MXXXXXXXXXXXXXXXXXXX18, S =>
                           MXXXXXXXXXXXXXXYFLXX, B => MXXXXXXXXXXXXXXXXXXX19, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXLL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX17 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX18 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXMXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXXXXXXX8 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX17 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXMXXXXX8, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLXXXXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX2, B => 
                           MXXXXXXXXXXXXXXYXX1, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXWXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL2, Y => 
                           MXXXXXXXXXXXXXXXXXXPXXLXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXXXXX2 : OR2 port map( A => MXMXXXX0, B =>
                           MXXXXXXXXXXXXXXXMXMXXXLXMXVXXXXFF, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXXXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXXXX5 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXX0 : NOR2A port map( A => MXMXXXXX(0), B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXXLXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXLX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXXLX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, C => MXXXXXXXXXXXXXXXJXMP
                           , Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX0 : NOR3 port map( A => XXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX7, C => MXXXXXXXXXXXXXXXXXXXX2, 
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX4 : OR2B port map( A => 
                           XXMXXXXX(6), B => MXXXXXXXXXXXXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXXXXXXX1 : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX5 : OR2B port map( A => 
                           XXMXXXXX(5), B => MXXXXXXXXXXXXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXXXXXXX2 : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX6 : OR2B port map( A => 
                           XXMXXXXX(4), B => MXXXXXXXXXXXXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXXXXXXX3 : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX7 : OR2B port map( A => 
                           XXMXXXXX(2), B => MXXXXXXXXXXXXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXXXXXXX4 : OR2B port map( A => 
                           MXMXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX8 : OR2B port map( A => 
                           XXMXXXXX(1), B => MXXXXXXXXXXXXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXXXXXXX5 : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX9 : OR2B port map( A => 
                           XXMXXXXX(0), B => MXXXXXXXXXXXXXXXXXXXPXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXXXXXXX6 : OR2B port map( A => 
                           MXMXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMXXFFHWX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXX8 : AO1A port map( A => MXXXXXXXXXXXXXXXXXXX17,
                           B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX00);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXFFXXXXXXXXXFXWXXX1 : NOR2A port map( A => 
                           XFXWX, B => MXXXXXXXXXXXXXXFXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXLXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXXLX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX, B => MXXXXXXXXXXXXXMXMPXXXXXXX,
                           Y => MXXXXXXXXXXXXXXXXXXMXMPXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL0, B => MXMXXXX0, Y
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL : OR2A port map( A => MXXXXXXXXXXXXXXYXX1
                           , B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXL2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXXXXXXX0 : NOR2A port map( A => MXMXXXX0, 
                           B => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXX3 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXPXXLXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXYXX1, B => MXXXXXXXXXXXXXXXXXXX21, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXYXXXXXX, B => MXXXXXXXXXXXXXXXXXXX21,
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXMMXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX1, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXMMX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXMMX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXMMX, C => 
                           MXXXXXXXXXXXXXXYXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXX1 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXYXXXXXX, C => MXXXXXXXXXXXXXXXXXXX21,
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXMXXXXXXXX0 : XAI1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX53, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXXXXXMXXXXXX : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXHXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXHXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXXX4 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => MXXXXXXXXXXXXXXXXXXXXXX
                           , Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXX2 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXHXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0, C => MXXXXXXXXXXXXXXYXX, 
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXXXXX4 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXHXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXHXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXHXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXXXXXXX1 : NOR2 port map( A => ramaddr(2), 
                           B => XXMXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXXXXXXX2 : NOR2B port map( A => XFXWX, B =>
                           ramaddr(2), Y => MXXXXXXXXXXXXXXXXXXFXWXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXXXXXXX10 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX00, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXMXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX9 : OR3B port map( A => XXMXXXXXXX,
                           B => MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, C => 
                           ramaddr(2), Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXL : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXL1, B => 
                           MXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXLXX2, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXLXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXL0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX10 : OR2B port map( A => 
                           XXMXXXXX(4), B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXXXXXXX3 : OA1B port map( C => 
                           MXXXXXXXXXXXXXMXMPXXXXX, A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXX : NOR2 port map( A => XXXXXPXXX, B
                           => MXXXXXXXXXXXXXXXXXXFXXXHX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX : NOR2 port map( A => XXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, B => 
                           MXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXMPXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX21 : MX2C port map( A => 
                           MXMXXXXXXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX22 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXWXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX42);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXXXXXXX10 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXMXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXX, C => MXXXXXXXXXXXXXXXXXX1, 
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPHWX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWXXX, B => 
                           MXXXXXXXXXXXXXXYXX, C => MXXXXXXXXXXXXXMXMPXXXXX, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPLWX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX11 : OR2B port map( A => 
                           XXMXXXXX(5), B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXXXXXXX12 : OR2B port map( A => 
                           XXMXXXXX(3), B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXXXMXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXMXXFFLWXXXXX, B => 
                           XXMXXXXX(0), Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXMXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXHX : DFN1P0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX6, CLK => 
                           XLXXPX, PRE => MXXXXXXXXXXXXXXXXXXXXX5, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXFXXXHXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXMXMXMXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX5, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXMXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFFXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX2, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXLXXX1, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMWX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXXXX, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => MXMWXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXX6, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX4, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXMXMXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXMXVXXXXFFXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXMXVXXXX, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXMXMPXXXX3, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXMXVXXXXFF);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXXXXXXX2, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => MXMXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX23 : DFN1E1C0 port map( D => XFXXXXXX(0),
                           E => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX24 : DFN1E1C0 port map( D => XFXXXXXX(1),
                           E => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWXXX1, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX25 : DFN1E1C0 port map( D => XFXXXXXX(2),
                           E => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX26 : DFN1E1C0 port map( D => XFXXXXXX(3),
                           E => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX27 : DFN1E1C0 port map( D => XFXXXXXX(4),
                           E => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX28 : DFN1E1C0 port map( D => XFXXXXXX(5),
                           E => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX29 : DFN1E1C0 port map( D => XFXXXXXX(6),
                           E => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX30 : DFN1E1C0 port map( D => XFXXXXXX(7),
                           E => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFXWX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXXXXXXX : DFN1E1C0 port map( D => 
                           MXMXXXXXXXXXXXXX1, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXMXXXXXXXXXXXXX2, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXMXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXMXXXXXXXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXXXXXXX3 : DFN1E1C0 port map( D => 
                           MXMXXXXXXXXXXXXX4, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXXXXXXX4 : DFN1E1C0 port map( D => 
                           MXMXXXXXXXXXXXXX0, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXXXXXXX5 : DFN1E1C0 port map( D => 
                           MXMXXXXXXXXXXXXX5, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXLXXXXXXXX6 : DFN1E1C0 port map( D => 
                           MXMXXXXXXXXXXXXX6, E => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXLWX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXLXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXPXLXXXXXX50);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX54, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXPXLXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX55, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXLXXXXXX00);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX56, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXLXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX57, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXLXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX58, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXLXXXXXX30);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX59, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXLXXXXXX40);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX60, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXLXXXXXX60);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX61, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXHXXXXXX40);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX62, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXHXXXXXX30);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX63, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXHXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX64, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXHXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX65, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXHXXXXXX60);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX66, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXPXHXXXXXX50);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX67, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX9, Q => 
                           MXXXXXXXXXXXXXPXHXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXPXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX7, CLK => XLXXPX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => 
                           MXXXXXXXXXXXXXPXHXXXXXX00);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2, 
                           CLK => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX9, Q => 
                           MXMXXXX1_0_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX8, CLK => XLXXPX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_1_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX9, CLK => XLXXPX, CLR 
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_2_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX10, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_3_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX11, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_4_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX12, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_5_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX13, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_6_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX14, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_7_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX15, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_8_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXX9 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX16, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXX1_9_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX17, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX10, Q => MXMXXXX1_10_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX18, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX10, Q => MXMXXXX1_11_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX19, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX10, Q => MXMXXXX1_12_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX20, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX10, Q => MXMXXXX1_13_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX21, CLK => XLXXPX, CLR
                           => MXXXXXXXXXXXXXXXXXXXXX10, Q => MXMXXXX1_14_port);
   MXXXXXXXXXXXXXXXMXMXXXLXMXMXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXX6, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXMXXXX1_15_port);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX1, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXXXXX2, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX6, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXVXXX5, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX1, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX3, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX2, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX4, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXX, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX9 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXX10 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX0, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX1, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX2, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX9 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX3, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXXXX10 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXXXXX4, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXFFXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX53, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX52, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX51, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX6 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX50, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX7 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX49, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX8 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX48, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX9 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX47, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX10 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX46, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX11 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX45, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX12 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX44, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX46, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX45, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX44, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX43, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX42, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX41, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX11 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX29, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX12 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX28, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX13 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX27, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX14 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX26, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX15 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX25, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX16 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX24, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX13, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX17 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX23, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX18 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX22, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX19 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX21, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXX20 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXX20, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX13 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX43, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX14 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX42, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX15 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX41, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX16 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX54, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX17 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX40, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXXXX18 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXXXX39, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXXX14, Q => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX15 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX16 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX13 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX14 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX5, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX15 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX16 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX17 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX18 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX7, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX19 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX7, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX20 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX28);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX21 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX29);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX22 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX27);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX23 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX23);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX30);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX25 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX7, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX24);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX26 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX31);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX27 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX10, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX25);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX28 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX5, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX32);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX29 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX6, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX26);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX30 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX11, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX31 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX32 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX33);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX33 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX34);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX34 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX0 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXX1, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX1 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX2 : AND3 port map( A => 
                           MXXXXXXXXXXXXXPXHXXXXXX60, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX50, C => 
                           MXXXXXXXXXXXXXPXHXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXX2, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX4 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX5 : AND2 port map( A => 
                           MXXXXXXXXXXXXXPXHXXXXXX60, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX50, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX6 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXX3, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX50, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX7 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX, C => 
                           MXXXXXXXXXXXXXPXHXXXXXX60, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX8 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXX2, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX60, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX9 : AND3 port map( A => 
                           MXXXXXXXXXXXXXPXHXXXXXX30, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX20, C => 
                           MXXXXXXXXXXXXXPXHXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX10 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXX4, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX49);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX11 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXPXHXXXXXX30, C => 
                           MXXXXXXXXXXXXXPXHXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX12 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX13 : AND3 port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX40, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX60, C => 
                           MXXXXXXXXXXXXXPXHXXXXXX40, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX14 : AND3 port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX10, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX20, C => 
                           MXXXXXXXXXXXXXPXLXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXXX15 : AND3 port map( A => 
                           MXXXXXXXXXXXXXPXLXXXXXX50, B => 
                           MXXXXXXXXXXXXXPXLXXXXXX7, C => 
                           MXXXXXXXXXXXXXPXLXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXFXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX17 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX18 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX7, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX19 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX20 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX21 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX22 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX6, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX23 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX5, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX36);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX43);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX25 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX44);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX26 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX42);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX27 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX38);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX28 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX45);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX29 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX9, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX39);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX30 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX46);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX31 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX40);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX32 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX7, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX33 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX8, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX41);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX34 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX37);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX35 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX35);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX36 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX47);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX37 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX48);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXXX38 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXXXXXXX35 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXPXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX8, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX9, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX10, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX1, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX1,
                           C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX11, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX9, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX50);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX12, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX53);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX1,
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX51);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX6 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXXX7 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXX : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXX0 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXHXXXXXXXXXXX3 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXHXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXPXXLXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX5 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX9, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX6 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX10, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX11, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX12, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX13, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX11, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX9, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX14, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX15, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX3 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX12, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX16, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX4 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX10, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX8, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX5 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX14, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0
                           , C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX6 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX12, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX,
                           C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX7 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX14, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX15, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX8 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX11, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX13, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX14, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX9 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX10, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX13, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX10 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX13, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX16, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX11 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX16, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX18, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX12 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX15, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX19, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX13 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX9, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX1, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX14 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX10, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX1
                           , C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX17, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX15 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX17, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX18, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX16 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX
                           , C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX14, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX17 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX11, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0
                           , C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX18 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX8, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX17, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX20, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX19 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX12, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX1
                           , C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX20 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX9, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX10, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX17, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX21 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX,
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX22 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX12, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX23 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX10, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX1
                           , Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX25 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXX0
                           , Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX26 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX13, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX27 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX8, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX28 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXX
                           , Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX29 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX7, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX30 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX11, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX31 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX8, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX9, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX32 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX13, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX33 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXX, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX34 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX35 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX41, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX36 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX37 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX44, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX38 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX40, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX39 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX40 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX43, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX41 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX42, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX42 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX43 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX45, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX44 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX45 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX46 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX39, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX47 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX48 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX49 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX50 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX51 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX40, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX52 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX53 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX54 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX44, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX55 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX41, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX56 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX57 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX43, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX58 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX39, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX59 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX60 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX61 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX62 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX42, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX63 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX64 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX65 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX39, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX66 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX67 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX3, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX68 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX43, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX69 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX70 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX42, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX71 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX72 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX41, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX40, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX44, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX3 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXVXXXXX4, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX4 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX45, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX7 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX13, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXXX8 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX15, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX16, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX73 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX18, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX19, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX74 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX21, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX17, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX75 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX22, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX23, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX76 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX24);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX77 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX25, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX26, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX78 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX20, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX14, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX27);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX79 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX22, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX2, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX80 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX25, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX3, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX81 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX27, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX4, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX82 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX15, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX16, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX5);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX83 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX16, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX6, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX7, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX84 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX15, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX21, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX6, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX85 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX19, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX9, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX10, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX86 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX26, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX3, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX12, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX87 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX23, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX2, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX14, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX88 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX17, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX15, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX8, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX89 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX20, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX11, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX90 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX17, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX16, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX91 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX19, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX20, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX17);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX92 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX15, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX93 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX21, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX15, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX94 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX22, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX23, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX95 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX14, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX11, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX17, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX96 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX24, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX5, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX97 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX18, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX9, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX98 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX19, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX2,
                           C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX18, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX99 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX13, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX18, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX19, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX100 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX18, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22, C 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX13, Y 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX101 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX55);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX102 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX7, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX25, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX62);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX103 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX18, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX63);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX104 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX8, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX61);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX105 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX9, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX57);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX106 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX26, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX64);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX107 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX10, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX14, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX58);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX108 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX65);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX109 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX11, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX21, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX59);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX110 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX21, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX66);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX111 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX12, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX17, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX60);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX112 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX13, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX19, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX56);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX113 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX14, B 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX2,
                           Y => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX54);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX114 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX22, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX67);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX115 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX24, Y 
                           => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX116 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX50, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX117 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX47, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX8);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX118 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX53, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX119 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX49, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX11);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX120 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX4);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX121 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX52, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX122 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX51, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX123 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX124 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX55, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX125 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX126 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX54, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX127 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX48, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX128 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX46, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX129 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX130 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX131 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX132 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX49, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX133 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX134 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX135 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX53, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX25);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX136 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX50, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX23);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX137 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX46, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX138 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX52, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX26);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX139 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX48, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX140 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX13);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX141 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX142 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXXX);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX143 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX54, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX144 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX51, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX22);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX145 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX47, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX146 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX147 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX48, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX7);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX148 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX54, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX18);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX149 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX150 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX46, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX10);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX151 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX52, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX12);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX152 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX153 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX51, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX2);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX154 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXXX155 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX50, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX14);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX5 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX6 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX49, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX6);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX7 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX53, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX3);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX8 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX47, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX9);
   MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXXX9 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXPXXXXXVXXXXX55, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXWXXXXXXXXXXXXXXMPXXXXX2);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity XYXX0001 is

   port( MXXXXXXXXXXXXXMXMXXXX, XLXXPX, MXXXXXXXXXXXXXXXXXXXXXX : in std_logic;
         MXXXXXXXXXXXXXXXXXXXXX, XXXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  XXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXXXXX0, XXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXX1, XXXXXXXX2
         , MXXXXXXXXXXXXXXXXXXXXX2 : out std_logic;  MXXXXXXXXXXXXXXXXXXXX, 
         MXMXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXX : out std_logic;
         MXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, MXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXWXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXXXXXXXWXXX : out std_logic;  MXXXXXXXXXXXXXXYXX, 
         MXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXX1
         , MXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXXXXXFXWXXXXX, XFXXXXXXXXXX, XFXXXXXXXXXX0, 
         MXXXXXXXXXXXXXMXMPXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXVXX, 
         MXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX1, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXX7, 
         MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX8, XFXXXXXXXXXXX, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXX11,
         MXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXX13, 
         MXXXXXXXXXXXXXMXMPXXXXXXX0, MXXXXXXXXXXXXXXXXXXX14, 
         MXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXX15, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXX16, 
         MXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXXXXXX19
         , MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXXXX7, 
         MXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXX20, 
         MXXXXXXXXXXXXXXXXXXXXXXVXX0, MXXXXXXXXXXXXXXYXXXX, 
         MXXXXXXXXXXXXXXXXXXX21 : in std_logic;  MXXXXXXXXXXXXXXXXXPXWXXXXWXXX 
         : out std_logic;  XFXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXFXXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXYXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4, 
         MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6 :
         out std_logic;  MXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXFXWXXX, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXX, MXXXXXXXXXXXXXXXXXXX23, 
         MXXXXXXXXXXXXXXXXXXPXXXXXXXX, MXXXXXXXXXXXXXXYXXXX1, 
         MXXXXXXXXXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXXXX25, MXXXXXXXXXXXXXXXXXXX26
         , MXXXXXXXXXXXXXXXXXXX27, MXXXXXXXXXXXXXXXXXXX28, 
         MXXXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXX29 : in std_logic;  
         MXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXX7, 
         MXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXX10 : 
         out std_logic;  MXXXXXXXXXXXXXXXXXXX30, MXXXXXXXXXXXXXXXXXXXXXXXVXX0, 
         MXXXXXXXXXXXXXXXXXX11, MXMXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXX12, 
         MXXXXXXXXXXXXXXXXXX13 : in std_logic;  MXXXXXXXXXXXXXXXXXX14 : out 
         std_logic;  MXMXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX1, 
         MXMXXXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXXXX3, MXMXXXXXXXXXXXXXXX4, 
         MXMXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXXYXXXX2, 
         MXXXXXXXXXXXXXMXMPXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXXXXXX32, MXXXXXXX : in std_logic;  
         MXXXXXXXXXXXXXXXXLXXXXXXX, MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX, 
         MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXX11, 
         MXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXVXX, 
         MXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXX33, 
         MXXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXXXX : in 
         std_logic;  MXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXX0, 
         MXXXXXXXXXXXXXXYFLXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX12 : in 
         std_logic;  MXMXXXXX : out std_logic_vector (7 downto 0);  
         MXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, 
         MXXXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXFXXXXXXXXXX0 : in std_logic; 
         MXXXXXXXXXXXXXXXMXXX : out std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXX1 : 
         in std_logic;  MXXXXXXXXXXXXXXXMXXX0, MXXXXXXXXXXXXXXXMXXX1, 
         MXXXXXXXXXXXXXXXMXXX2 : out std_logic;  MXMXXXXXXXXXXXXXXX6, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, MXMXXXXXXXXXXXXXXX7, 
         MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX9, MXMXXXXXXXXXXXXXXX10, 
         MXXXXXXXXXXXXXXXXXXX34, MXXXXXXXXXXXXXXXXXXX35, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXXXXXXXX14, 
         MXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2, 
         MXXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXXXX15 : in std_logic;
         MXXXXXXXXXXXXXXXXLXXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXXX36, 
         MXXXXXXXXXXXXXXXXXXX37, MXMXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXXXX16
         , MXXXXXXXXXXXXXXXXXXXXXXXVXX2, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, 
         MXXXXXXXXXXXXXXXXXXX38, MXXXXXXXXXXXXXXXXXXX39, MXXXXXXXXXXXXXXXXXXX40
         , MXXXXXXXXXXXXXXXXXXXXXXXVXX3, MXXXXXXXXXXXXXXXXXXXX5, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX2 : in std_logic;  MXXXXXXXXXXXXXXXMXXX3 : 
         out std_logic;  XFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX3, 
         MXXXXXXXXXXXXXXFXXXXXXXXXX4 : in std_logic;  ramaddr : in 
         std_logic_vector (5 downto 0);  MXXXXXXXXXXXXXXXMXXX4, 
         MXXXXXXXXXXXXXXXMXXX5 : out std_logic;  MXXXXXXXXXXXXXXYXXXXXX, 
         MXXXXXXXXXXXXXMXMPXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXX2, 
         MXXXXXXXXXXXXXXYXX0 : in std_logic;  MXXXXXXXXXXXXXXXXXVXXXXXX, 
         MXXXXXXXXXXXXXXXXXXXXXXWXXX0, MXXXXXXXXXXXXXXXXXXXXXXWXXX1, 
         MXXXXXXXXXXXXXXXMXXX6, MXXXXXXXXXXXXXXXJXMP, MXXXXXXXXXXXXXXXXVXLXX : 
         out std_logic;  MXXXXXXXXXXXXXXXXXXXX6, MXMXXXXXXXXXXXXX0, 
         MXMXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX7, 
         MXXXXXXXXXXXXXXFXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXX8, 
         MXXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXXX10 : in std_logic;  
         MXXXXXXXXXXXXXXXXLXXXXXXX1 : out std_logic;  MXXXXXXXXXXXXXXXXXXXX11 :
         in std_logic;  MXXXXXXXXXXXXXXXXLXXXXXXX2 : out std_logic;  
         MXXXXXXXXXXXXXXXXXXXX12, 
         MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX : in std_logic);

end XYXX0001;

architecture SYN_USE_DEFA_ARCH_NAME of XYXX0001 is

signal MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWX, 
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXLXXXXXXXX, XXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX0, XXXXXXXX00, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX1, MXXXXXXXXXXXXXXXXXXXXX00, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX2, XXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX3, MXXXXXXXXXXXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX4, XXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX5, MXXXXXXXXXXXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX, MXXXXXXXXXXXXXXXXLXXXYFLXXXX, 
   MXXXXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX7, MXXXXXXXXXXXXXXXXLXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX9, MXXXXXXXXXXXXXXXXLXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX10, MXXXXXXXXXXXXXXXXLXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX, 
   MXXXXXXXXXXXXXXXXXXXXXXWXXX2, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXMXXXXX, MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXX19, MXXXXXXXXXXXXXXXXLXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXXXXX21, MXXXXXXXXXXXXXXXXLXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX, MXXXXXXXXXXXXXXXXLXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXXX1,
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXX0
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX0, MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX0,
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX, MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXX,
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX79, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX, MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXM, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX, MXXXXXXXXXXXXXXXXLXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX1
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX3
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXLXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX7, MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXXXX0
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXX, MXXXXXXXXXXXXXXXXLXXPXWXXX2, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX4, MXXXXXXXXXXXXXXXXLXXPXWXXX3, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX6
   , MXXXXXXXXXXXXXXXXLXXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXXMXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXX23, MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXMXXX, MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX2,
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2
   , MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX5, MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX6, MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX0
   , MXXXXXXXXXXXXXXXXLXXXXXMXXX0, MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXXMXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX4, MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX7,
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX5, MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX8,
   MXXXXXXXXXXXXXXXXLXXXXXXXX9, MXXXXXXXXXXXXXXXXLXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXMXXX2, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX10, MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX6
   , MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX13, MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX1,
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX1, MXXXXXXXXXXXXXXXXLXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXMXXX3, MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXX, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX3,
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX10, MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXMXXX4, MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX8, MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX14
   , MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX16, MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX3, MXXXXXXXXXXXXXXXXLXXXXXMXXX5, 
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX7, MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXXXVXXXXXXX, MXXXXXXXXXXXXXXXXLXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXXMXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX1, MXXXXXXXXXXXXXXXXLXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXMXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXX, MXXXXXXXXXXXXXXXXLXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX2, MXXXXXXXXXXXXXXXXLXXMXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXMXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX3, MXXXXXXXXXXXXXXXXLXXMXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX12
   , MXXXXXXXXXXXXXXXXLXXXXMXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX4, MXXXXXXXXXXXXXXXXLXXMXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX14, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX15
   , MXXXXXXXXXXXXXXXXLXXXXMXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXX, MXXXXXXXXXXXXXXXXLXXMXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX17, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX18
   , MXXXXXXXXXXXXXXXXLXXXXMXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXM, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX2, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX3, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXX24, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX7, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX8, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX8, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX13, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX4,
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXX25, 
   MXXXXXXXXXXXXXXXXLXXXXXXVXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXVXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX14, MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXX, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX14
   , MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX18, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX6,
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX7, MXXXXXXXXXXXXXXXXLXXMXXXMXXX, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX, MXXXXXXXXXXXXXXXXLXXMXXXMXXX0, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX0, MXXXXXXXXXXXXXXXXLXXMXXXMXXX1, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX1, MXXXXXXXXXXXXXXXXLXXMXXXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX2, MXXXXXXXXXXXXXXXXLXXMXXXMXXX3, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX3, MXXXXXXXXXXXXXXXXLXXMXXXMXXX4, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX,
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX7, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX9, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXX26, 
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXX27, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX2, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX21, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX11, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX23, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX8,
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX24, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX25, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX26, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX27, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX28, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX9,
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXMXXX, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX29
   , MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX14, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX30, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX31, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX10
   , MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX32, 
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX11, MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX12, MXXXXXXXXXXXXXXXXLXXMXXXMXXX5, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, MXXXXXXXXXXXXXXXXLXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX15, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX16, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX17, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX18, MXXXXXXXXXXXXXXXXLXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX1, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX9,
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX14, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX3, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX12
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX5, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX15
   , MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXMXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXX28, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX16, MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX1, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX19, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX20, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX8
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX21
   , MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX22, MXXXXXXXXXXXXXXXXLXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX9, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX23
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX10, MXXXXXXXXXXXXXXXXLXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX11, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX3
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXX7, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX24, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX25, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX26, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX14, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX33, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX19, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX34, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX35, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX36, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX37, 
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXLXXXPXXXMXXX0, 
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX14, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXMXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX16, MXXXXXXXXXXXXXXXXLXXXXXXX29, 
   MXXXXXXXXXXXXXXXXLXXXXXXX30, MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX17, MXXXXXXXXXXXXXXXXLXXXXXXX31, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXX32, 
   MXXXXXXXXXXXXXXXXLXXXXXXX33, MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX18, MXXXXXXXXXXXXXXXXLXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXX34, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXX35, 
   MXXXXXXXXXXXXXXXXLXXXXXXX36, MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXX37, MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXX38, MXXXXXXXXXXXXXXXXLXXXXXXX39, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXX40, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX0, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX1, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX2, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX3, MXXXXXXXXXXXXXXXXLXXXXMXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXMXXX8, MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX0, MXXXXXXXXXXXXXXXXLXXXXMXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXMXXX10, MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX2, MXXXXXXXXXXXXXXXXLXXXXMXXX11, 
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXMXXX12, MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX3, MXXXXXXXXXXXXXXXXLXXMXXXMXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX8, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX6, MXXXXXXXXXXXXXXXXLXXMXXXMXXX7, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX1
   , MXXXXXXXXXXXXXXXXLXXXXXXXXVXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXMXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXX41, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX0, MXXXXXXXXXXXXXXXXLXXMXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXX42, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXX43, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXX44, MXXXXXXXXXXXXXXXXLXXXXXXX45, 
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXX46, 
   MXXXXXXXXXXXXXXXXLXXXXXXX47, MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXX48, MXXXXXXXXXXXXXXXXLXXXXXXX49, 
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXX50, 
   MXXXXXXXXXXXXXXXXLXXXXXXX51, MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXX52, MXXXXXXXXXXXXXXXXLXXXXXXX53, 
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXX54, 
   MXXXXXXXXXXXXXXXXLXXXXXXX55, MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXX56, MXXXXXXXXXXXXXXXXLXXXXXXX57, 
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX7, MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX8
   , MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXX, MXXXXXXXXXXXXXXXXXPXWXXXXWXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXX0, MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXXXXX
   , MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX3, MXXXXXXXXXXXXXXXXLXXPXWXMXXX, 
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX0, MXXXXXXXXXXXXXXXXLXXPXWXMXXX0, 
   MXXXXXXXXXXXXXXXXLXXPXWXMXXX1, MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX2, MXXXXXXXXXXXXXXXXLXXPXWXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXPXWXMXXX3, MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX0, MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX2, MXXXXXXXXXXXXXXXXLXXPXXXXYXXXX, 
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX18, MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX20, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX3, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX1, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX21, MXXXXXXXXXXXXXXXXLXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX3, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX20, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXXXX0, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX21, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX15, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX7,
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX5, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX0, MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX0, MXXXXXXXXXXXXXXXXLXXMXXXMXXX8, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX1, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX2, MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXMXXX13, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXMXXX14, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX24, MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX25, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX37, MXXXXXXXXXXXXXXXXLXXXXXXX58, 
   MXXXXXXXXXXXXXXXXLXXXXXXX59, MXXXXXXXXXXXXXXXXLXXXXXXX60, 
   MXXXXXXXXXXXXXXXXLXXXXXXX61, MXXXXXXXXXXXXXXXXLXXXXXXX62, 
   MXXXXXXXXXXXXXXXXLXXXXXXX63, MXXXXXXXXXXXXXXXXLXXXXXXX64, 
   MXXXXXXXXXXXXXXXXLXXXXXXX65, MXXXXXXXXXXXXXXXXLXXXXXXX66, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXLXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXX67, MXXXXXXXXXXXXXXXXLXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX27, MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX28, MXXXXXXXXXXXXXXXXLXXXXXXXX29, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXXX30, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX31, MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX32, MXXXXXXXXXXXXXXXXLXXXXXXXX33, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXLXXXXXXXX34, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX35, MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXLXXXXXXXX36, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX37, MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX38, MXXXXXXXXXXXXXXXXLXXXXXXXX39, 
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXLXXXXXXXX40, 
   MXXXXXXXXXXXXXXXXLXXMXXXMXXX9, MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXMXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX15, MXXXXXXXXXXXXXXXXLXXXXXXX68, 
   MXXXXXXXXXXXXXXXXLXXXXXXX69, MXXXXXXXXXXXXXXXXLXXXXXXX70, 
   MXXXXXXXXXXXXXXXXLXXXXXXX71, MXXXXXXXXXXXXXXXXLXXXXXXX72, 
   MXXXXXXXXXXXXXXXXLXXXXXXX73, MXXXXXXXXXXXXXXXXLXXXXXXX74, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXLXXXXXXXXMXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX10, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX11
   , MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX12, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXVXXXXXX, MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXLXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, 
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXX, MXXXXXXXXXXXXXXXXLXXXXXXX75, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX41, MXXXXXXXXXXXXXXXXLXXXXXXXX42, 
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXX76, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, 
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXX77, 
   MXXXXXXXXXXXXXXXXLXXXXXXX78, MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, MXXXXXXXXXXXXXXXXLXXMXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXX1, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXMXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX39, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXLXXMXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXXXMXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXX79, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX, MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX5, MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX0, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX7, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX1, MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX7, MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX9, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX3, MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX9, MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX11, MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX5, MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXX0, 
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX11, MXXXXXXXXXXXXXXXXLXXXXMXMXXX, 
   MXXXXXXXXXXXXXXXXLXXXXMXMXXX0, MXXXXXXXXXXXXXXXXLXXXXMXMXXX1, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX43, MXXXXXXXXXXXXXXXXLXXXXMXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXMXMXXX3, MXXXXXXXXXXXXXXXXLXXXXMXMXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX, MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXXX00, 
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX2, MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXYFLXX0, MXMXXXXX0_1_port, MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX, 
   MXMXXXXX0_0_port, MXMXXXXX0_2_port, MXXXXXXXXXXXXXXXXLXXMXXXXX13, 
   MXMXXXXX0_6_port, MXMXXXXX0_7_port, MXXXXXXXXXXXXXXXXLXXXXVXXXX0, 
   MXMXXXXX0_5_port, MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXLXXXXXXXX44, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX5, MXXXXXXXXXXXXXXXXLXXXXXXXX45, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX46, MXXXXXXXXXXXXXXXXLXXXXXXXX47, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX48, MXXXXXXXXXXXXXXXXLXXXXXXXX49, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX50, MXXXXXXXXXXXXXXXXLXXXXXXXX51, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX52, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX39, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX21, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX11, MXXXXXXXXXXXXXXXXLXXXXXXXX53, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX23, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX12, MXXXXXXXXXXXXXXXXLXXXXXXXX54, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX25, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX27, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX28, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX13, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX29, MXXXXXXXXXXXXXXXXLXXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX15, MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX7, MXXXXXXXXXXXXXXXXLXXXXXXXX55, 
   MXXXXXXXXXXXXXXXXLXXXXMXXX15, MXXXXXXXXXXXXXXXXLXXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX17, MXXXXXXXXXXXXXXXXLXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX19, MXXXXXXXXXXXXXXXXLXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX21, MXXXXXXXXXXXXXXXXLXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXXXX7, MXXXXXXXXXXXXXXXXLXXPXWXXX4, 
   MXXXXXXXXXXXXXXXXLXXPXWXXX5, MXXXXXXXXXXXXXXXXLXXPXWXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX40, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX41
   , MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX42, 
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX43, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX44
   , MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX45
   , MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX46, MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX3,
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX4, MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX10, MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX12, MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX14, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX19
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX25, MXXXXXXXXXXXXXXXXLXXXXXXX80, 
   MXMXXXXX0_3_port, MXMXXXXX0_4_port, MXXXXXXXXXXXXXXXXLXXMXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXXXXX81, MXXXXXXXXXXXXXXXXLXXXXXXX82, 
   MXXXXXXXXXXXXXXXXLXXXXXXX83, MXXXXXXXXXXXXXXXXLXXXXXXX00, 
   MXXXXXXXXXXXXXXXXLXXXXXXX85, MXXXXXXXXXXXXXXXXLXXXXXXX86, 
   MXXXXXXXXXXXXXXXXLXXXXXXX87, MXXXXXXXXXXXXXXXXLXXXXXXX88, 
   MXXXXXXXXXXXXXXXXLXXXXXXX89, MXXXXXXXXXXXXXXXXLXXXXXXX90, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXXXXXX56, MXXXXXXXXXXXXXXXXLXXXXXXX91, 
   MXXXXXXXXXXXXXXXXLXXXXXXX92, MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX27, MXXXXXXXXXXXXXXXXLXXXXXXX93, 
   MXXXXXXXXXXXXXXXXLXXXXXXX94, MXXXXXXXXXXXXXXXXLXXXXXXX95, 
   MXXXXXXXXXXXXXXXXLXXXXXXX96, MXXXXXXXXXXXXXXXXLXXXXXXX97, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXX16, MXXXXXXXXXXXXXXXXLXXXXXXX98, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, MXXXXXXXXXXXXXXXXXXXXXXWXXX00, 
   MXXXXXXXXXXXXXXXXXXXXXXWXXX10, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX40, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX41, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX42, MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX43
   , MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX31, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX44, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX45, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX21, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX9, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX10, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX24, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX32, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX26, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX27, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX25, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX26, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX27, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX28, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX29, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX30, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX31, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX28, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX29, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX30, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX5, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX17, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX24, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX18, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX19, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX32, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX33, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX34, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX35, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX36, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX37, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX38, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX39, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX40, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX41, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX42, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX2, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX21, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX43, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX31, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX32, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX33, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX34, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX35, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX36, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX37, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX6, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX11, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX12, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX0, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX13, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX14, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX7, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX22, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX25, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX44, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX3, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX23, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX45, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX38, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX1, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX39, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX8, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX15, 
   MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX16 : std_logic;

begin
   MXXXXXXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXXXX17;
   XXXXXXXX <= XXXXXXXX3;
   XXXXXXXX0 <= XXXXXXXX00;
   MXXXXXXXXXXXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXXXXXXXX00;
   XXXXXXXX1 <= XXXXXXXX10;
   MXXXXXXXXXXXXXXXXXXXXX1 <= MXXXXXXXXXXXXXXXXXXXXX18;
   XXXXXXXX2 <= XXXXXXXX20;
   MXXXXXXXXXXXXXXXXXXXXX2 <= MXXXXXXXXXXXXXXXXXXXXX20;
   MXXXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXX15;
   MXXXXXXXXXXXXXXXXXXXXXXWXXX <= MXXXXXXXXXXXXXXXXXXXXXXWXXX2;
   MXXXXXXXXXXXXXXXXXPXWXXXXWXXX <= MXXXXXXXXXXXXXXXXXPXWXXXXWXXX0;
   MXXXXXXXXXXXXXXXXLXXXXXXX <= MXXXXXXXXXXXXXXXXLXXXXXXX78;
   MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX0;
   MXXXXXXXXXXXXXXXXXXXXXXXX <= MXXXXXXXXXXXXXXXXXXXXXXXX1;
   MXXXXXXXXXXXXXXXXXXXXXXXX0 <= MXXXXXXXXXXXXXXXXXXXXXXXX00;
   MXXXXXXXXXXXXXXYFLXX <= MXXXXXXXXXXXXXXYFLXX0;
   MXMXXXXX <= ( MXMXXXXX0_7_port, MXMXXXXX0_6_port, MXMXXXXX0_5_port, 
      MXMXXXXX0_4_port, MXMXXXXX0_3_port, MXMXXXXX0_2_port, MXMXXXXX0_1_port, 
      MXMXXXXX0_0_port );
   MXXXXXXXXXXXXXXXXLXXXXXXX0 <= MXXXXXXXXXXXXXXXXLXXXXXXX00;
   MXXXXXXXXXXXXXXXXXXXXXXWXXX0 <= MXXXXXXXXXXXXXXXXXXXXXXWXXX00;
   MXXXXXXXXXXXXXXXXXXXXXXWXXX1 <= MXXXXXXXXXXXXXXXXXXXXXXWXXX10;
   
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXMXMXXXXXXXXXXXXXXX : OR2 port map( A 
                           => MXXXXXXXXXXXXXMXMXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX, Q => XXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX0, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX0, Q => XXXXXXXX00);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX2 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX3 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX0, Q => XXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX4 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX5 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX0, Q => XXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX6 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXPXWXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXLXXXYFLXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXMXXXXXXXXXXXXX, E => MXXXXXXXXXXXXXXXXXX15, CLK =>
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => MXXXXXXXXXXXXXXXXXXX0, C 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX0 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => XXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => XXXXXXXX00, Y =>
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => XXXXXXXX10, Y =>
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX5 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => XXXXXXXX20, Y =>
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX6 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX13, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX7 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX14, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX8 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX15, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX9 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX16, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX10 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX17, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX11 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX18, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXMXMXXXXXXXXXXXXX : OR2 port map( A =>
                           MXXXXXXXXXXXXXMXMXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXMXMXXXXXXXXXXXXX0 : OR2 port map( A 
                           => MXXXXXXXXXXXXXMXMXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXFXWXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXPXXXXXXVXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYXX, B => MXXXXXXXXXXXXXXXXXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXYXXXPXXXXMXXXVXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX1, B => MXXXXXXXXXXXXXXXXXXXXX4
                           , Y => MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXYXXXPXXXXXXXXXYXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX1, B => MXXXXXXXXXXXXXXXXXXXXX4
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, B 
                           => MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, B
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX1 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, 
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXPXXXXXXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX3, B => MXXXXXXXXXXXXXXXXXXXX1, 
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXXXXXXX0 : AND2 port map( A => XFXXXXXXXXXX
                           , B => XFXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX79, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXM, B => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX4 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXYFLXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX79, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX5 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXXXX, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX6 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXXXXXXX7 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXFXXXXXXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX1 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX4 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX5 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX4 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXFXXXXXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX5 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX6 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX6 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX10 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX11 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX12 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX13 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX7 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX9 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX10 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX14 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX15 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX16 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXXXXXXX17 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX6, B => MXXXXXXXXXXXXXXXXXXX7, C
                           => MXXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXXXXXX5,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX7, Y
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX5, B => MXXXXXXXXXXXXXXXXXXX6,
                           C => MXXXXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX0 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXXXVXXXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXXXVXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           XFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX7 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX8 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX10 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX11 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX12 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX13 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX14 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX15 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX16 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX17 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX18 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXXXXXXX19 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXM, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX2 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX5 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX6 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX7 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX8 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX9 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX10 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX11 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX12 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX13 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXXXXXXX2 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX14 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX15 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX16 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX17 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX18 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXXXXXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXXXXXXXMXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXXXXXXXMXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXXXXXXXMXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXXXXXXXMXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX19 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX20 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX21 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX22 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX13, B => MXXXXXXXXXXXXXXXXXXX10,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX23 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX24 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX25 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX27, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX26 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX26);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX27 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX27);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX28 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX28);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX29 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX29, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX30);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX30 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX31, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX29);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX31 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX32);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX32 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX31);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX, B
                           => MXXXXXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX4 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX,
                           B => MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX6 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX7 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX8 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX9 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX10 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX11 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX12 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0
                           , B => MXXXXXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX13 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1
                           , B => MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX13);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX14 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX15 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX16 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX17 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX18 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX19 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX20 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX21 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX22 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX23 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2
                           , B => MXXXXXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX26);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXXXXXXX24 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3
                           , B => MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX33 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX33, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX19, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX34);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX34 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX36, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX33);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX35 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX37);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX36 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX35);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXX37 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXYFLXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXMXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX36);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX : AXOI5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX29, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXXXX : AXOI5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX31, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXXXX0 : AXOI5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX32, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXXXX1 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX33, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXXXX2 : AXOI5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX34, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXXXX3 : AXOI5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX35, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXXXX4 : AXOI5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXXXX5 : AXOI5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXXXX6 : AXOI5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX40, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXXXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXXXXXXX1 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXXXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXXXXXXX4 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXXXXXXX5 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXXXX2 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXXXX3 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX3 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXXXXXVXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXVXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXXXXXVXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXXXXXVXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXXXXXVXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXXXX0 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXXXX1 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX42, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXXXX2 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX43, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX44, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX45, Y => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXXXX0 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX46, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX47, Y => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXXXX1 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX48, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX49, Y => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXXXX2 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX50, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX51, Y => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXXXX3 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX52, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX53, Y => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXXXX4 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX54, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX55, Y => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXXXX5 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX56, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX57, Y => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : AO1A port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX3 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX4 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX5 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX6 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX7 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX8 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXXXXXXXX : OR2A port map( A 
                           => MXXXXXXXXXXXXXXYXXXX, B => MXXXXXXXXXXXXXXXXXXX21
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXX, B => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXXXXXXX0 : NOR3 port map( A => 
                           XFXXXXXXXXXX1, B => XFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX0, B => MXXXXXXXXXXXXXXYXX, Y =>
                           MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX3);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXLXXXVXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXLXXXVXXXXX0 : OA1A port map( A => XXXXXXXX00, B 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXLXXXVXXXXX1 : OA1A port map( A => XXXXXXXX3, B 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX0, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXLXXXVXXXXX2 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX1, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXLXXXVXXXXX3 : OA1A port map( A => XXXXXXXX20, B 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX1, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXLXXXVXXXXX4 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXLXXXVXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX00, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX2, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXLXXXVXXXXX6 : OA1A port map( A => XXXXXXXX10, B 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX3, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, B => XFXXXXXXXXXX, C => 
                           XFXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX);
   MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXXXXXXX : XOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX17, B => XXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXXXXXXX0 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX00, B => XXXXXXXX00, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX);
   MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX18, B => XXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX20, B => XXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXXXXX : XOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXXXXX2 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXXXXX3 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXXXXX4 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX5 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX6 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX26, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX7 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXMXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4
                           , C => MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX20, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXX5 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX21, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXX6 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX1);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXX2 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX2);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXYFLXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX1 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX5, B => MXXXXXXXXXXXXXXXXXXX22
                           , C => MXXXXXXXXXXXXXXXXLXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX, C => 
                           MXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXXXVXXXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX2 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3A port map( 
                           A => MXXXXXXXXXXXXXXYXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX24, C => MXXXXXXXXXXXXXXXXXXX25,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXXXXXXXXXXXXXXXXX : OR3B port map( A 
                           => MXXXXXXXXXXXXXXYXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX26, C => MXXXXXXXXXXXXXXXXXXX25,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX37);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX26);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX58, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX59, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX60);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX61, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX62, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX63);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX1 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX64, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX65, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX66);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX3 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX27, B => MXXXXXXXXXXXXXXXXXXX28,
                           C => MXXXXXXXXXXXXXMXMPXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX3 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0,
                           C => MXXXXXXXXXXXXXXXXXXXXXXVXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX28, B => MXXXXXXXXXXXXXXXXXXX27,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXX9, C => MXXXXXXXXXXXXXXXXXXX29
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXX67);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX27, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX0 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX28, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX29, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX1 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX31, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX2 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX32, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX33, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX3 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX34, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX35, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX4 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX5 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX39, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXXXVXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXXXVXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXXXVXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX11 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX7, A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX68, Y => 
                           MXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXX0 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX6, A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX69, Y => 
                           MXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXX1 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX5, A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX70, Y => 
                           MXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXX2 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX4, A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX71, Y => 
                           MXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXX3 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX3, A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX72, Y => 
                           MXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXX4 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX2, A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX73, Y => 
                           MXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX74);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXXXXXX0 : NOR2A port map( A 
                           => MXXXXXXXXXXXXXXXXXXX30, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXX8 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXVXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX27);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXX0 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXX1 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXX3 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXX4 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXX5 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX12);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXX3 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX3);
   MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXX1 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXVXXXXX7, A => 
                           MXXXXXXXXXXXXXXXXLXXXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXX : OR3B port map( 
                           A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXYXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXX0 : OR3 port map( 
                           A => MXXXXXXXXXXXXXXXXLXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX1 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXPXWXVXXXXXXMXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXYFLXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXPXWXVXXXXXXMXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXYFLXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX75, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX18, C =>
                           MXXXXXXXXXXXXXXXXLXXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX42);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, B => 
                           MXMXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXV : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXVXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXX);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXX1 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX39, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXX2 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXXXX3 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXX5 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX1, A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX76, Y => 
                           MXXXXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, B => 
                           MXMXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, B => 
                           MXMXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXX1 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, B => 
                           MXMXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXX2 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, B => 
                           MXMXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, B => 
                           MXMXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXX1 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, B => 
                           MXMXXXXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXFXWXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXX5 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXVXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX31, B => MXXXXXXXXXXXXXXYXXXX2, 
                           C => MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX26, C => 
                           MXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX2, B => MXXXXXXXXXXXXXXXXXXX32, 
                           C => MXXXXXXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX77);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXXXVXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX0 : NOR2B port map( A => MXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXX78, Y => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXXXXXXXX0 : OR2B port map( A 
                           => MXXXXXXXXXXXXXXYXXXX2, B => MXXXXXXXXXXXXXXXXXXX7
                           , Y => MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXXXXXVXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXVXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXXXXXX1 : NOR2 port map( A =>
                           MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => MXXXXXXXXXXXXXXXXXXXXX3, 
                           C => MXXXXXXXXXXXXXXXXXXXXXXXVXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXVXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXX0 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX18, A => 
                           MXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX33, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX2 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX79);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXX : NOR2 port map( A 
                           => MXXXXXXXXXXXXXXXXLXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXX1 : AO1D port map(
                           A => MXXXXXXXXXXXXXXXXLXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXX3 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXVXXXX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX33, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXX2 : OR2B port map(
                           A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXX3 : OR2 port map( 
                           A => MXXXXXXXXXXXXXXXXLXXXYFLXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX11, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXX);
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXXXXXXX10 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX39);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX5 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX12, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXMXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX13, S => 
                           MXXXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX79, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX4);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXXXX0 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX5);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXXXX1 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX6);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXXXX2 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX7);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXXXX3 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX8);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX9);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXXXX5 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX10);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXXXX6 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX0);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX1);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX2);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX2 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX3);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX3 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX4);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX4 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX9);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXM);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX6);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX7);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXXXXXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX4 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX8);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXXXXXXX1 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX5 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX9);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXXXXXXX2 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX6 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX10);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXXXXXXX3 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX7 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX11);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXXXXXXX4 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXX0);
   MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXXXXXXX5 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXXVXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXXXXX : MX2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXXXXYXXXX, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXX4);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXX : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX1, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX1, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX00, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXX2 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXX3 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXPXWXVXXXXXXMXXX1 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXYFLXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXMXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXM);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX5 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXX : OR2A port map( A => MXMXXXXX0_1_port,
                           B => MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX12, B => MXMXXXXX0_0_port, C 
                           => MXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX4);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX6 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXX0 : OR2A port map( A => MXMXXXXX0_2_port
                           , B => MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX12, B => MXMXXXXX0_1_port, C 
                           => MXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX6);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX7 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX7);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX8 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXX1 : OR2A port map( A => MXMXXXXX0_6_port
                           , B => MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX6);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX2 : OR2A port map( A => 
                           MXMXXXXX0_7_port, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX3 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX12, B => MXMXXXXX0_6_port, C 
                           => MXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX8 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXMXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXMXX);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXXMXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXFXXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX1 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXMXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX5);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXFXXXXXXXMXXXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXFXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX2 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXMXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX3 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX3 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXX0 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX5 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXX1 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXXMXXXXXXXX2 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX4 : OR3A port map( A => 
                           MXMXXXXX0_5_port, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX5 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXMXXXXXXXX3 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX5 : OR3A port map( A => 
                           MXMXXXXX0_6_port, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX7 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX6);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXX2 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXMXXXXXXXX4 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX6 : OR3A port map( A => 
                           MXMXXXXX0_7_port, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX9 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX1 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX12);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX2 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXX : AO1 port map( A => MXXXXXXXXXXXXXXXXXXX13, B
                           => MXXXXXXXXXXXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX : XAI1 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXXXXXXX : XAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX15);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXX18, B => MXXXXXXXXXXXXXXXXXXX19,
                           C => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX0 : XAI1 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX17, C => 
                           MXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX0 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXX18, B => MXXXXXXXXXXXXXXXXXXX19,
                           C => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX1 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX1 : XAI1 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX2 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXX18, B => MXXXXXXXXXXXXXXXXXXX19,
                           C => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX2 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, C => 
                           MXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX2 : XAI1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, C => 
                           MXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX9);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX4 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXX18, B => MXXXXXXXXXXXXXXXXXXX19,
                           C => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX5 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX3 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX3 : XAI1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX10, C => 
                           MXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX7);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX6 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX18, B => MXXXXXXXXXXXXXXXXXXX19,
                           C => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX7 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX4 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX8 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX18, B => MXXXXXXXXXXXXXXXXXXX19,
                           C => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX9 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX10 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX5 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX4 : XAI1 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, C => 
                           MXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX6);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX11 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX18, B => MXXXXXXXXXXXXXXXXXXX19,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYFLXX0, B => MXXXXXXXXXXXXXXXXXXX13, 
                           Y => MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX12 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXMXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX44, B => 
                           MXXXXXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX5 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX4, B
                           => MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX15);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX6 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX16);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX45, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX46, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX47, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX48, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX49, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX50, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX51, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXX5 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX52, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX3 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX13);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX4 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX5 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX9);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX6 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX53, B => 
                           MXXXXXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX7 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX7);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX8 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX54, B => 
                           MXXXXXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX9 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX10 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX11 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXMXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX12 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX13 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX14 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXMXXX15 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXXXXXXX3 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX7 : OR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX6, B
                           => MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX17);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX8 : OR2B port 
                           map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXMXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX55, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXXXX4 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXXXX5 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXXXX6 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX2, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX14);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX3, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX13);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX4, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX7);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX5, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX8);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX1, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX9);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX5 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX10);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX6 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX11);
   MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXXXXXXX13 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXMXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX1 : AX1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX2 : AXO5 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXMXXX : OR3C port map( A => MXXXXXXXXXXXXXXFXXXXXXXXXX0
                           , B => XFXXXXXXXXXX, C => MXXXXXXXXXXXXXXXXLXXXXXX0,
                           Y => MXXXXXXXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX4, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXX0 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXX, Y => MXXXXXXXXXXXXXXXMXXX0
                           );
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX5, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXX2 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX2);
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX00, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX3);
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX6, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX39);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXX0 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX40);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX41);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX42);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXX3 : MX2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX43);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXX4 : MX2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX44);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXX5 : MX2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX45);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXX6 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, S => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX46);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX : MX2B port map( A => MXMXXXXXXXXXXXXXXX6, S
                           => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX0 : MX2B port map( A => MXMXXXXXXXXXXXXXXX7, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX1 : MX2B port map( A => MXMXXXXXXXXXXXXXXX8, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX2 : MX2B port map( A => MXMXXXXXXXXXXXXXXX9, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX3 : MX2B port map( A => MXMXXXXXXXXXXXXXXX2, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX4 : MX2B port map( A => MXMXXXXXXXXXXXXXXX1, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX5 : MX2B port map( A => MXMXXXXXXXXXXXXXXX10,
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX6 : MX2B port map( A => MXMXXXXXXXXXXXXXXX8, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXX0, B => 
                           MXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX7 : MX2B port map( A => MXMXXXXXXXXXXXXXXX9, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXX0, B => 
                           MXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX8 : MX2B port map( A => MXMXXXXXXXXXXXXXXX2, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXX0, B => 
                           MXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX9 : MX2B port map( A => MXMXXXXXXXXXXXXXXX1, 
                           S => MXXXXXXXXXXXXXXXXXXXXXXXVXX0, B => 
                           MXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXX10 : MX2B port map( A => MXMXXXXXXXXXXXXXXX10
                           , S => MXXXXXXXXXXXXXXXXXXXXXXXVXX0, B => 
                           MXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX9 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXVXXXX : AX1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXVXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX6 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXXXXXPXWXVXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX33, C => MXXXXXXXXXXXXXXXXXXX31,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXPXWXVXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXPXXXXXXXXXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX2, B => MXXXXXXXXXXXXXXXXXXX34, 
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX10 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXWXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX, B => MXXXXXXXXXXXXXXXXXXX35, Y
                           => MXXXXXXXXXXXXXXXXLXXXXXXX80);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXX3, Y => MXXXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXX : NOR2 port map( A => 
                           MXMXXXXX0_3_port, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX64);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX4 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX65);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX5 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXX3, C => MXMXXXXX0_2_port, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX41);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXX0 : NOR2 port map( A => 
                           MXMXXXXX0_4_port, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX61);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX6 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX62);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX7 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXX4, C => MXMXXXXX0_3_port, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX42);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX58);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX8 : NOR2 port map( A => 
                           MXMXXXXX0_5_port, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX59);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX9 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXX4, C => MXMXXXXX0_4_port, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX43);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX10 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX79);
   MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXVXXXXXXXXXX11 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX28);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXYXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXYXXXPXXXXXXXXXYXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXYXXXPXXXXMXXXVXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX : AO1B port map( A => 
                           MXXXXXXXXXXXXXXYXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX1, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX81, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXX : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX83, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX47);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX00, B => 
                           MXXXXXXXXXXXXXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX78);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXX1 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX85, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX49);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXX2 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX86, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX51);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXX3 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX87, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX53);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXX4 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX88, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX55);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXX5 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX89, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX57);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXX : AX1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX37, B => 
                           MXXXXXXXXXXXXXXXXXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXXXXVXXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX40);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX29, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX90, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX38);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX39);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX0 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX31, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX36);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX67, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX30, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX37);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX32, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX90, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX3 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX34);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX4 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX67, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX33, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX35);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX5 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX90, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX32);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX6 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX33);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX7 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX30);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX8 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX67, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX31);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX9 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX90, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX28);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX10 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX29);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX11 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX40, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX26);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX12 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX67, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX27);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX12 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX13 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX75, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXXXX0, C 
                           => MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX41);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX14 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX15 : NOR2A port map( A => 
                           MXMXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX56);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXPXXXXXXVXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXYXX, B => MXXXXXXXXXXXXXXXXXXX4, Y =>
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXYXXXPXXXXXXVXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYXX, B => MXXXXXXXXXXXXXXXXXXXXX14, Y
                           => MXXXXXXXXXXXXXXXXLXXXXVXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX67, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX3 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX13 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXX7 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX15);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, B => MXMXXXXX0_0_port
                           , Y => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX0 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX7, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => MXMXXXXX0_1_port,
                           Y => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX1 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX8, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => MXMXXXXX0_2_port,
                           Y => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX2 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX9, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => MXMXXXXX0_3_port,
                           Y => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX10, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => MXMXXXXX0_4_port,
                           Y => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => MXMXXXXX0_5_port,
                           Y => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX5 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX12, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => MXMXXXXX0_6_port,
                           Y => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX6 : MX2C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX13, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, B => MXMXXXXX0_7_port,
                           Y => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX7 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX91, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX8 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX14, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX9 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX15, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX10 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX16, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX11 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX92, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX12 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX17, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX13 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX18, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXX14 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX93, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX : MX2B port map( A => MXMXXXXXXXXXXXXXXX11
                           , S => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX94);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX0 : MX2B port map( A => MXMXXXXXXXXXXXXXXX6
                           , S => MXXXXXXXXXXXXXXXXXXXXXXXVXX0, B => 
                           MXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX95);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX1 : MX2B port map( A => 
                           MXMXXXXXXXXXXXXXXX11, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX0, B => 
                           MXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX96);
   MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX2 : MX2B port map( A => MXMXXXXXXXXXXXXXXX7
                           , S => MXXXXXXXXXXXXXXXXXXXXXXXVXX0, B => 
                           MXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX97);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX4 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXX38, B => MXXXXXXXXXXXXXXXXXXX20,
                           C => MXXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXX : AX1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX90);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXMXXXX : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX0, S => MXXXXXXXXXXXXXXXXXXXXX15,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX31);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXMXXXX0 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX2, S => MXXXXXXXXXXXXXXXXXXX39, B
                           => MXXXXXXXXXXXXXXXXLXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX34);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXMXXXX1 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX3, S => MXXXXXXXXXXXXXXXXXXX39, B
                           => MXXXXXXXXXXXXXXXXLXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX37);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXMXXXX2 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX12, S => MXXXXXXXXXXXXXXXXXXX39, 
                           B => MXXXXXXXXXXXXXXXXLXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX40);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXMXXXX : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX11, S => MXXXXXXXXXXXXXXXXXXX39, 
                           B => MXXXXXXXXXXXXXXXXLXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX29);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXMXXXX3 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX1, S => MXXXXXXXXXXXXXXXXXXX39, B
                           => MXXXXXXXXXXXXXXXXLXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX32);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXMXXXX4 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX13, S => MXXXXXXXXXXXXXXXXXXX39, 
                           B => MXXXXXXXXXXXXXXXXLXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX35);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXMXXXX5 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX4, S => MXXXXXXXXXXXXXXXXXXX39, B
                           => MXXXXXXXXXXXXXXXXLXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX38);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX16 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX56, A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX75);
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXXXX14 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX38, B => MXXXXXXXXXXXXXXXXXXX40,
                           C => MXXXXXXXXXXXXXXYFLXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXX3 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX81);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX5 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX30);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX6 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX33);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX7 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX36);
   MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXXX8 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX39);
   MXXXXXXXXXXXXXXXXLXXXXMXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXX9 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXMXXXXXXXX4 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXMXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXPXXXXPXWXVXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXYFLXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXVXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXXXX17 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXXXVXXXXXXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2, B => 
                           XFXXXXXXXXXXX0, C => MXXXXXXXXXXXXXXXXLXXXXXXXX42, Y
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX7);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX7 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXXXXX6 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX37, B => MXXXXXXXXXXXXXXXXXXX39,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXX98, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX45);
   MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXXXXXXX3 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX8 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXXXXXXX9 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXMXXX8);
   MXXXXXXXXXXXXXXXXLXXMXXXMXXXXXXXXXX8 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXMXXXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXXXXXXX7 : OR3A port map( A => 
                           MXMXXXXX0_4_port, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXMXXXXXXXX5 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXX4 : OR3C port map( A => ramaddr(4), B => 
                           ramaddr(5), C => MXXXXXXXXXXXXXXXXLXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX2, B => ramaddr(5), Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXX5 : OR3C port map( A => ramaddr(4), B => 
                           ramaddr(5), C => MXXXXXXXXXXXXXXXXLXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXXLXXPXWXMXXXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYFLXX0, B => ramaddr(5), Y => 
                           MXXXXXXXXXXXXXXXXLXXPXWXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => MXXXXXXXXXXXXXXXXXXX0, C 
                           => MXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXMXMPXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXYXXXXXX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXXXXXXXXX : OR2A port map( A 
                           => MXXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXYXX0, Y => MXXXXXXXXXXXXXXXXXVXXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXX4 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX00, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXX5 : NOR2 port map( A => ramaddr(3), B 
                           => ramaddr(2), Y => MXXXXXXXXXXXXXXXXXXXXXXWXXX00);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXXXXXXX6 : NOR2 port map( A => ramaddr(1), B 
                           => ramaddr(0), Y => MXXXXXXXXXXXXXXXXXXXXXXWXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX7 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXLXXXXMXXX6 : OR3C port map( A => ramaddr(4), B => 
                           ramaddr(5), C => MXXXXXXXXXXXXXXXXLXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXXXXXXX10 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXVXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXMXXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXMXMXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXMXMXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXVXXXXXXXXX : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX77, A => 
                           MXXXXXXXXXXXXXXXXXXX32, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXVXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXXXXXXX2 : AO1A port map( A => 
                           MXXXXXXXXXXXXXMXMXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXPXXXXXXXXMXMXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXMXMXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXWX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXX);
   MXXXXXXXXXXXXXXXXLXXXXJXMPXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXLXXXXXXXX, CLK => XLXXPX
                           , CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXJXMP);
   MXXXXXXXXXXXXXXXXLXXXXXVXLXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXMXFXXXXXXMXX, E => 
                           MXXXXXXXXXXXXXXYXX0, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX0, Q => MXXXXXXXXXXXXXXXXVXLXX)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX95, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX91);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX96, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX97, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX2 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX10, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX3 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX11, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX92);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX4 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX12, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX5 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX13, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX6 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX14, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX80, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX93);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX7 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX8 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX94, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX9 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX10 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX11 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX12 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX7, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX13 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX14 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXYXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX82, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           MXMXXXXXXXXXXXXX, E => MXXXXXXXXXXXXXXXXXX15, CLK =>
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXMXXXXXXXXXXXXX0, E => MXXXXXXXXXXXXXXXXXX15, CLK 
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX2 : DFN1E0C0 port map( D => 
                           MXMXXXXXXXXXXXXX1, E => MXXXXXXXXXXXXXXXXXX15, CLK 
                           => XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXPXWXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXX4, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX4);
   MXXXXXXXXXXXXXXXXLXXPXWXXXXXXXX0 : DFN1E1C0 port map( D => XFXXXXXXXXXXX0, E
                           => MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXX6, Q => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX5);
   MXXXXXXXXXXXXXXXXLXXPXWXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX0, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX3);
   MXXXXXXXXXXXXXXXXLXXPXWXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXPXWXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX00);
   MXXXXXXXXXXXXXXXXLXXPXWXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXPXWXXXXWX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX6);
   MXXXXXXXXXXXXXXXXLXXPXWXXXXXXXX3 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX3, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXX2);
   MXXXXXXXXXXXXXXXXLXXPXWXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXPXWXXXYXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXYFLXX0);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX2);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX3);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX4);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX7, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX5);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX1);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX4 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX7, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX6);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX5 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX10, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX7);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX6 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX11, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX0 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX1 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX2 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX8, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX3 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX4 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX5 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX0, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX6 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXYXXXXX, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXWXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX7 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXXXX, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXMXXXXX0_0_port);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX8 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXX, Q => 
                           MXMXXXXX0_1_port);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX9 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX0, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXXX0_2_port
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX10 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXXX0_3_port
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX11 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXXX0_4_port
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX12 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXXX0_5_port
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX13 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXXX0_6_port
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXX14 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXYXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXMXMXXXXXXX, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX9, Q => MXMXXXXX0_7_port
                           );
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX7 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX3, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX12, CLK => XLXXPX, CLR =>
                           MXXXXXXXXXXXXXXXXXXXX9, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX10);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX8 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX2, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX74, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX9, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX8);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX9 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX1, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX74, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX9);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX10 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX66, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX74, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX11 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX63, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX74, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX13);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX12 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX60, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX74, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX0);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX13 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX0, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX74, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX14);
   MXXXXXXXXXXXXXXXXLXXMXXXXXXXXXX14 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXXYXXXXX, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX74, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX15 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX7, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX80, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX73);
   MXXXXXXXXXXXXXXXXLXXXXXXX3 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX6, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX80, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX16 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX80, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX76);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX17 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX10, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX80, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX72);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX18 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX80, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX71);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX19 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX5, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX80, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX70);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX20 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX4, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX80, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX69);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX21 : DFN1E0C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX11, E => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX80, CLK => XLXXPX, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX68);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX22 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX3, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX46);
   MXXXXXXXXXXXXXXXXLXXXXXXX4 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX15, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX10, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX00);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX23 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX1, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX44);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX24 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX0, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX48);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX25 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX14, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX50);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX26 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX13, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX52);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX27 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX12, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX54);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX28 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXXX2, CLK => XLXXPX, 
                           CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX56);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX29 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXX7, CLK => XLXXPX,
                           CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX83);
   MXXXXXXXXXXXXXXXXLXXXXXXX5 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX13, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX30 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX12, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX98);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX31 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX11, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX85);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX32 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX10, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX86);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX33 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX9, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX11, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX87);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX34 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX8, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX88);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXX35 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXXLXXXXXXXXXXXXX7, CLK => 
                           XLXXPX, CLR => MXXXXXXXXXXXXXXXXXXXX12, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX89);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX8 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX6 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX,
                           B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, 
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2, 
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX7 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX0, 
                           B => MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX1, C
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3, 
                           Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX8 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0, 
                           B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX1, 
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX9 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1, 
                           B => MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX1, Y
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX10 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX11 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX9 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX10 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX11 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX12 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX13 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX14 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX12 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX13 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, 
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX,
                           Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX14 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX1
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, 
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX15 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2
                           , B => MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX2,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX1
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX16 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX5, 
                           Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX0
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX17 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX7
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX4, 
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX18 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2, 
                           B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX1,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX19 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX8
                           , B => MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX2,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX20 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX21 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX22 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX8
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX23 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX7
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX0
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX15 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX2
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX16 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX17 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX18 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX1
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX19 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX20 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX25 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX26 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX53);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX27 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX0,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX54);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX28 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX29 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX30 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3
                           , B => MXXXXXXXXXXXXXXYFLXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX2
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX21 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX3
                           , B => MXXXXXXXXXXXXXXYFLXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX31 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX0, 
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX32 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX, 
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX33 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX34 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX1
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX22 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX4
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX5
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX6
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX7
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX8
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX8
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX3 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX5
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6, 
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX7, 
                           Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX2
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX4 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXX1, 
                           B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, 
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX9, 
                           Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX5 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX4
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, 
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6, 
                           Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX6 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX7
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX10,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX11,
                           Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX3
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX7 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX4
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX8 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX6
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, C
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX10,
                           Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX9 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX8
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX2
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX3
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX10 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX9
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX39, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX5
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX11 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX4
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX6
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX7
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX12 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, 
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX2
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX13 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX3
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX7
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX14 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX15 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX9
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX2,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX16 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3, 
                           B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX55);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX17 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX10, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX12,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX18 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4, 
                           B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX0, Y
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX19 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX11, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX20 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5, 
                           B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX21 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6, 
                           B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX8, 
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX22 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX42, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX9
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX23 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX46, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX25 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX44, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX26 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX45, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX27 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX28 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX41, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX29 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX41, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX30 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX45, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX6
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX31 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX42, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX32 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX9
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX33 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX44, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX5
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX34 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX4
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX35 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX46, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX7
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX36 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX45, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX10)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX37 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX41, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX4
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX38 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX44, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX46, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX11)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX43, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX42, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX6
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXPXXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX5
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX23 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX4
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX35 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX25 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX44);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX36 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX37 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX5
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX, Y
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX6 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX7 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX0
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX38 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX6
                           , B => MXXXXXXXXXXXXXXXXLXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX40, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX13,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX40, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX0 : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX41, B 
                           => MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX2,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX13)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX1 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX13,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX40, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX2 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX3,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX42, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX3 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX2, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX4 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX43, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX31, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX5 : OR3A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX31, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX43, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX6 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX43, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX31, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX7 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX44);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX8 : NOR3A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX45);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX9 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX39 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX4, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX40 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX6, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX7, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX41 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX5, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX8, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX42 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX9, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX10, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX43 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX9, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX14,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX8
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX44 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX6, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX9
                           , Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX45 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX10, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX46 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX7, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX9
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX11, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX47 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX5, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX13, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX48 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX4, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX10, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX14, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX49 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX10, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX15, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX50 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX10, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX8
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX16, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX51 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX8, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX13, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX12, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX52 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX12, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX16,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX18, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX14)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX53 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX11, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX14,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX17, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX54 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX12, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX1, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX52);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX55 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX13, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX15,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX49);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX56 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX14, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXX45);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX57 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX15, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX5,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX51);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX58 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX16, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX16,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX46);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX59 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX17, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX14,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX47);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX60 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX18, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX2, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXX50);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX61 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX19, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX4,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXX48);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX62 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX63 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX64 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX65 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX66 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX67 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX68 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX69 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX70 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX71 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX72 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX73 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX74 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX75 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX76 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX77 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX78 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX26 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX20, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX9
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX27 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX28 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX29 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX30 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXVXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX8
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX31 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX16)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX32 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX33 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXX0);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX34 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXMXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX11 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX17,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX45, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX12 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX44, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX13 : OR3A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX44, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX17)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX14 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX44, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX10 : NOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX11 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX13, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX18,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX19, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX19)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX12 : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX13 : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX18,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX14 : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX20,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX18)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX15 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX18,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX16 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX6,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX17 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX19,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX31, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX18 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX20,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX19 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXYFLXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX20 : OR3A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXYFLXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX19, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX20)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX21 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXYFLXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX22 : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX40, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX40, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX7)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX23 : AO1A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX41, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX8,
                           C => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX24 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX21,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX40, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX25 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX7,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX42, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX26 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX8,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX27 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX43, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX28 : OR3A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX43, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX8)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX29 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX43, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX15 : XNOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX9,
                           B => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX45, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX16 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX44, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX17 : OR3A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX44, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX9)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX18 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX44, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX30 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX11, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX20, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX31 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX14, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX10
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX21, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX32 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX20, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX22,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX33 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX21, B 
                           => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX34 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX22, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX10
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX35 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX36 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX37 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX39, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX38 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX39 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX40 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX41 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX42 : OR3 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX9, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX10
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX43 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX15, 
                           B => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX44 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX39, B 
                           => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX9);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX45 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX39, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX46 : AOI1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX11
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX12, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX22, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX42);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX47 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX12
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX23, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX11
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX48 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX23, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX11
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX40);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX49 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX24, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX12
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX41);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX50 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX43);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX51 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX52 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX53 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX54 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX55 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX56 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX57 : OR3 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX12
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX58 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX59 : AND2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX13, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX14, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX60 : AOI1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX13
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX15, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX24, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX32);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX61 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX14, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX25, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX26, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX62 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX13, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX13
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX25, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX14
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX63 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX0, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX15
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX27, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX13
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX64 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX25, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX13
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX65 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX26, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX14
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX66 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX27, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX15
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX67 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX26);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX68 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX69 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX70 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX27);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX71 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX72 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX73 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX74 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX75 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX76 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX77 : OR3A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX15
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX78 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX79 : AND2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX15, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX16, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX80 : AOI1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX16, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX28, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX31);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX81 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX16, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX29, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX30, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX82 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX15, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX29, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX17
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX83 : AO1 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX1, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX18
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX31, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX84 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX28, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX16
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX85 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX29, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX17
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX86 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX30, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX18
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX87 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX9, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX29);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX88 : XOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX89 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX28);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX90 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX30);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX91 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX92 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX93 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX94 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX95 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX15, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX31);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX96 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX29);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX97 : OR3A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX18
                           );
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXXXXXXXXXXX98 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX17, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX18, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX20, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX21, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX19, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX22, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX23, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX24, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX3 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX23, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX19
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX32, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX33);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX4 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX20, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX34, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX5 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX17, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX35, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX6 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX21, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX34, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX36, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX37);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX7 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX19, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX38, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX8 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX18, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX35, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX39, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX38);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX9 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX17, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23,
                           C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX40, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX10 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX24, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX32, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX41, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX42);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX11 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX22, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX38, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX37, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX40);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX12 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX2, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX21
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX43, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX19
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX13 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXX18, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX19
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX42, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX14 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX31, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX15 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX32, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXX23,
                           Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX16 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX
                           , B => MXXXXXXXXXXXXXXXXLXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX17 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX33, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX20
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX18 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX34, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX21
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX19 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX35, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX19
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX20 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX36, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXXX4, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX21 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX37, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX33, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX22 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX35);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX23 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX31);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX24 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX25 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX34);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX26 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX36);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX27 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX33);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX28 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX37);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX29 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX32);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX30 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX31 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX32 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX33 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX34 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX35 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX36 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX37 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX36);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXXX38 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX39);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX20, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX34);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX35);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX1 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX41);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX2 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX43);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX3 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX32);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX4 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX21
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX5 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX12);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX6 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXXLXXMXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX11);
   MXXXXXXXXXXXXXXXXLXXXXXXMXXXXXXXXXX7 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX25, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX19 : XOR2 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX20 : XNOR2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX21 : NOR3 port 
                           map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX7, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXLXXXXXVXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX22 : AND2 port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX13);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX23 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX14);
   MXXXXXXXXXXXXXXXXLXXXXMXXXXXXXXXLXXXXXLXXPXXXXXXXXLXXXXXVXXX24 : NOR2A port 
                           map( A => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX0 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX22
                           , B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX25, C 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX44, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX1 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX3, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX23
                           , C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX45, Y 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX22
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX2 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX38, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX22
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX3 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX1, B 
                           => MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX4 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX39, B 
                           => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX23
                           , Y => MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX5 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX6 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX39);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX7 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXLXXXMXXXXX38);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX8 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX9 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXPXXXXXXXYXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX10 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX45);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX11 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX27, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXXX44);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX12 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX15, C => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXXXXXXYXXXXXXXX23
                           );
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX13 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX32, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX16);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX14 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXX15);
   MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX15 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXPXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX32, Y => 
                           MXXXXXXXXXXXXXXXXLXXXWXXXXXXXXXXXXXXMPXXXXXX8);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,PROASIC3;

use IEEE.std_logic_1164.all;
use PROASIC3.components.all;

entity CORE8051 is
generic (
USE_OCI     : integer := 0;
USE_UJTAG   : integer := 0;
TRACE_DEPTH : integer := 0;
TRIG_NUM    : integer := 0;
NRSTOUT     : integer := 0;
EN_FF_OPTS  : integer := 0
);

   port( port0i, port1i, port2i, port3i : in std_logic_vector (7 downto 0);  
         port0o, port1o, port2o, port3o : out std_logic_vector (7 downto 0);  
         memdatai : in std_logic_vector (7 downto 0);  memdatao : out 
         std_logic_vector (7 downto 0);  memaddr : out std_logic_vector (15 
         downto 0);  ramdatai : in std_logic_vector (7 downto 0);  ramdatao, 
         ramaddr : out std_logic_vector (7 downto 0);  sfrdatai : in 
         std_logic_vector (7 downto 0);  sfrdatao : out std_logic_vector (7 
         downto 0);  sfraddr : out std_logic_vector (6 downto 0);  membank : in
         std_logic_vector (3 downto 0);  TraceA : out std_logic_vector (7 
         downto 0);  TraceDI : out std_logic_vector (19 downto 0);  TraceDO : 
         in std_logic_vector (19 downto 0);  nreset, clk, clkcpu, clkper, int0,
         int1, int0a, int1a, int2, int3, int4, int5, int6, int7, rxd0i, t0, t1 
         : in std_logic;  nrsto, nrsto_nc, clkcpu_en, clkper_en, movx, rxd0o, 
         txd0 : out std_logic;  mempsacki, memacki : in std_logic;  mempsacko, 
         mempsrd, memwr, memrd, ramwe, ramoe, sfrwe, sfroe : out std_logic;  
         TCK, TMS, TDI : in std_logic;  TDO : out std_logic;  TRSTB, BreakIn : 
         in std_logic;  BreakOut, dbgmempswr, TrigOut, AuxOut, TraceWr : out 
         std_logic);

end CORE8051;

architecture SYN_verilog of CORE8051 is

   component XYXX0008
      port( XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0 : in std_logic;  
            XXXXXXXXXXXXXXXXXJXXXXX : out std_logic;  XLX, XXXXXXXX : in 
            std_logic;  JXXXXX, XXXXXX : out std_logic;  
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX : in std_logic;  XXXXXXXX0 
            : out std_logic;  MXMXXXXXXXX : in std_logic;  MXMXXXX : in 
            std_logic_vector (15 downto 0);  XXXXXXX : in std_logic_vector (19 
            downto 0);  XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXPX, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, XXXXXXXX1, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXP, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH : in std_logic;  MXMXXXX0 
            : in std_logic_vector (3 downto 0);  MXMXXXXXXXX0, XXXXXXXX2, 
            MXMXXXXXXXX1, MXMXXXXXXXX2, XXXXXXXX3, XXXXXXXX4, XXXXXXXX5 : in 
            std_logic;  XXXXXXXXP : out std_logic;  
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX1, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX2, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX3, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX4, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX5, 
            XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX6, XXXXXX0 : in 
            std_logic;  XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, 
            XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, 
            XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1, 
            XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2, 
            XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3, 
            XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4, 
            XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5, 
            XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6 : out std_logic;  
            XXXXXXXX6, XXXXXXXX7 : in std_logic;  XXXXXPXWX, XXXXXPXXX, 
            XXXXXXXX8 : out std_logic;  XXXXXXX0, XXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXXXXXX, MXMPXXXXX : in std_logic);
   end component;
   
   component XYXX0007
      port( XLXXPX, MXXXXXXXXXXXXXXXXXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXXX0 : out 
            std_logic;  MXMXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXPXXXXXX, MXXXXXXXXXXXXXXXXXXFXXXHX : out 
            std_logic;  MXXXXXXXXXXXXXXXXXFXXXHXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX 
            : in std_logic;  MXXXXXXXXXXXXXXYXLXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  
            MXXXXXXXXXXXXXXYXLXXXXXX0, MXXXXXXXXXXXXXXYXLXXXXXX1 : out 
            std_logic;  MXXXXXXXXXXXXXXXXPPMX, MXXXXXXXXXXXXXXXXXXMXMPXXXX : in
            std_logic;  MXXXXXXXXXXXXXXYXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXXXXX7, 
            MXXXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXXXX11 : out 
            std_logic;  MXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  
            MXXXXXXXXXXXXXXMWXXXXXXX, MXXXXXXXXXXXXXXMWXXXXXXX0 : out std_logic
            ;  MXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXLLXX, MXXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXYXXXX, MXXXXXXXXXXXXXXYXXXX0
            , MXXXXXXXXXXXXXXYXXXX1, MXXXXXXXXXXXXXXXXXFXXXHX, 
            MXXXXXXXXXXXXXXYXLXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXPXXXXXX
            , MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, MXMXXXXXXXXXXXXXXX0, 
            MXMXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXMXMPXXXX, MXXXXXXXXXXXXXXXXXXXMXMPXXXX0, 
            MXXXXXXXXXXXXXXXXXXXPXXXXXX0, MXMXXXXXXXXXXXXXXX2, 
            MXMXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXMXMPXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0 : out std_logic;  
            MXMXXXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXXXX6, 
            MXMXXXXXXXXXXXXXXX7, MXMXXXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXXPXXXXXX1, MXMXXXXXXXXXXXXXXX8, 
            MXMXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXX0, XXXXXXXXXXXXXXXXXX : in
            std_logic;  MXVX : out std_logic;  MXMXXXXXXXXXXXXXXX10, 
            MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, MXMXXXXXXXXXXXXXXX11, 
            MXMXXXXXXXXXXXXXXX12, MXMXXXXXXXXXXXXXXX13 : in std_logic;  
            MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX : out std_logic;  
            MXMXXXXXXXXXXXXXXX14, MXMXXXXXXXXXXXXXXX15 : in std_logic;  
            MXXXXXXXXXXXXXXYXLXXXX0, MXXXXXXXXXXXXXXYXX : out std_logic;  
            MXMXXXXXXXXXXXXXXX16, MXMXXXXXXXXXXXXXXX17 : in std_logic;  
            MXXXXXXXXXXXXXXYXLXXXX1, MXXXXXXXXXXXXXXYXLXXXX2, 
            MXXXXXXXXXXXXXXYXX0, MXXXXXXXXXXXXXXYXXXX2, MXXXXXXXXXXXXXXYXX1 : 
            out std_logic;  MXMXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXMXMPXXXXXXX0, 
            MXXXXXXXXXXXXXMXMPXXXXXXX1 : in std_logic;  
            MXXXXXXXXXXXXXXXXYXLXXXXX : out std_logic;  MXMXXXXXXXXXXXXXXX19, 
            MXMXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXXXPXXLXX, 
            MXXXXXXXXXXXXXXXXXMXVXWXXX, MXXXXXXXXXXXXXXXXXXX1 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXLL : out std_logic;  XXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXXXPFF, MXMXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXX0,
            MXMXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXX3, 
            MXMXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXX6 : in 
            std_logic;  MXXXXXXXXXXXXXXXXXX1 : out std_logic;  
            MXXXXXXXXXXXXXMXMPXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXMXMXXXLXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXMWXXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX : 
            in std_logic;  MXXXXXXXXXXXXXXXXYXLXXXXX0, 
            MXXXXXXXXXXXXXXXXYXLXXXXX1, MXXXXXXXXXXXXXXXXYXLXXXXX2, 
            MXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXXXX2 : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX3 :
            in std_logic;  MXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXXX7, 
            MXXXXXXXXXXXXXXXXXXXXX8 : out std_logic);
   end component;
   
   component XYXX0006
      port( MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, XLXPXX, MXXXXXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXFXWXXX, XFXXXXXXXXXX,
            MXXXXXXXXXXXXXXXXXPXWXXXXWXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXX0 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXXVXX : in std_logic;  MXXXXXXXXXXXXXXXXXXXXX
            : out std_logic;  MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, 
            MXXXXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXXXX0 : out
            std_logic;  MXXXXXXXXXXXXXXYXXXX, MXXXXXXXXXXXXXXYXXXX0 : in 
            std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9, MXXXXXXXXXXXXXXXXPXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12, MXXXXXXXXXXXXXXXXVXXXXXX, 
            MXXXXXXXXXXXXXXXXVXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXFX, 
            MXXXXXXXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXXXVXXXXXX1, 
            MXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXX0 : out std_logic;  
            MXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXL : out 
            std_logic;  MXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXFX0 : in 
            std_logic;  MXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXVXXXXXX2, 
            MXXXXXXXXXXXXXXXXVXXXXXX3, MXXXXXXXXXXXXXXXXXX1 : out std_logic;  
            MXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXX2 : in 
            std_logic;  MXXXXXXXXXXXXXXXXXXFXXXXX, MXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXPXXXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXFXWXXX
            : in std_logic;  MXXXXXXXXXXXXXXXXXXX2 : out std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXXXPXXXXXXXX1, MXXXXXXXXXXXXXXXXPXXXXXXXX2 : out 
            std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXX2, 
            XXMXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXX4 : out std_logic;  
            XXXXX, MXXXXXXXXXXXXXXXXXXXXX2, XXXXX0, XXXX, XXXX0, XXXX1, XXXX2, 
            XXXX3, XXXX4, MXXXXXXXXXXXXXXXXXXXXX3 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXX4 : out std_logic;  
            MXXXXXXXXXXXXXXXXXFXXXHXXX, MXXXXXXXXXXXXXXXXXFXXXHX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX1 : in std_logic;  XFXXXXXX : in 
            std_logic_vector (7 downto 0);  XFXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXX4, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXXXXXXXX6 : in std_logic);
   end component;
   
   component XYXX0005
      port( MXXXXXXXXXXXXXXYXLXXXXXX, MXXXXXXXXXXXXXXYXLXXXXXX0 : in std_logic;
            MXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXXX3 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXFXXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0
            , MXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1, MXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXFXWXXXXX, MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX : 
            in std_logic;  MXXXXXXXXXXXXXXXXXXFXWXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXFXWXXX, XFXXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX0 : in 
            std_logic;  MXXXXXXXXXXXXXXXXXXFXWXXX0 : out std_logic;  XXXX : in 
            std_logic;  MXXXXXXXXXXXXXXXX1 : out std_logic;  XXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX4 : in std_logic;
            MXXXXXXXXXXXXXXXX2 : out std_logic;  MXXXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXYXLXXXXXX1, MXXXXXXXXXXXXXXYXLXXXX : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXMXXX : out std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
            XFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXX 
            : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXWXXX, 
            MXXXXXXXXXXXXXXLXXXVXX, MXXXXXXXXXXXXXXFXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXFXWXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXX3 : in 
            std_logic;  MXXXXXXXXXXXXXXFXXXXXXXMXXX0 : out std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXX, XFXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXXXXXXX7, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX8, MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX10, MXXXXXXXXXXXXXXFXXXXXXXXXXX11, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXXXXXXFXWXXX0 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXMXXX, MXXXXXXXXXXXXXXXXXXMXXXXX, 
            MXXXXXXXXXXXXXXXXXXMXXX0 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXFXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXX1 : out std_logic;  XFXWX : in std_logic;  
            MXXXXXXXXXXXXXXFX : out std_logic;  MXXXXXXXXXXXXXXXXXXXX6 : in 
            std_logic;  MXXXXXXXXXXXXXXFX0 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXX7 : in std_logic;  MXXXXXXXXXXXXXXXXVXX : out 
            std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXX6, 
            MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, XXMXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXMXXX1 : out std_logic;  XXMXXXXXXX0, XXMXXXXXXX1
            , XLXPXX, MXXXXXXXXXXXXXXXXXXXXXXX, XX, XX0, MXXXXXXXXXXXXXXXXXXXXX
            : in std_logic;  XFXXXXXX : in std_logic_vector (8 downto 2);  
            MXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXXXX3 : in std_logic);
   end component;
   
   component XYXX0004
      port( XLXPXX, MXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX : in 
            std_logic;  MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXXXXXXLXX, MXXXXXXXXXXXXXXLXXXVXX, 
            MXXXXXXXXXXXXXXXXXXXXX, XFXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX, 
            XFXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXLXXXXXXXXXX, MXXXXXXXXXXXXXXFXWXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX0 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXFXWXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXWXXX, MXXXXXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXX0 : out std_logic;  XFXXXXXXXXXX1, XXMXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXX, XFXXXXXXXXXXX, 
            XFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX5, MXXXXXXXXXXXXXXFXXXXXXXXXXX6, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX7, MXXXXXXXXXXXXXXFXXXXXXXXXXX8, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX9 : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXXX4 : out 
            std_logic;  MXXXXXXXXXXXXXXXXXXFXWXXX0, 
            MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, XFXWX, MXXXXXXXXXXXXXXXXVXX, 
            XXMXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX1 : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXXXX5, MXXXXXXXXXXXXXXFXXXXXXXXXXXX6 : out 
            std_logic;  MXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXMXX, 
            MXXXXXXXXXXXXXXLXXXVX, MXXXXXXXXXXXXXXLXXXVX0, 
            MXXXXXXXXXXXXXXXXXXXXXXXXX, XXXXX, MXXXXXXXXXXXXXXXXXXXXX0 : in 
            std_logic;  XXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX1 : in 
            std_logic;  XXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXX4, 
            MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXX6, 
            MXXXXXXXXXXXXXXXXXXXXX7 : in std_logic);
   end component;
   
   component XYXX0003
      port( MXXXXXXXXXXXXXXXXXXXXXX, XLXXPX, MXXXXXXXXXXXXXXXXXXXXXXXXX : in 
            std_logic;  XFXXXXXXXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX
            : in std_logic;  XFXXXXXXXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXMXMPXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXPXXXXXX : out 
            std_logic;  MXXXXXXXXXXXXXXXXXXXPXXXXXX0 : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXXX : out std_logic;  MXMXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX : out std_logic;  
            MXMXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXXXXXXPXXXXXX1 : 
            out std_logic;  MXXXXXXXXXXXXXMXMPXXXXXXX, MXMXXXXXXXXXXXXXXXXX, 
            MXMXXXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXX0, 
            MXMXXXXXXXXXXXXX1, MXMXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXX4, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX5, XFXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXXXXXX7, 
            XFXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXX8, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX9, XFXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXX 
            : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX2 : out std_logic;  MXXXXXXXXXXXXXXXXXX0
            : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX4 : out std_logic;  MXXXXXXXXXXXXXXXXXX1
            : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX6 : out std_logic;  MXXXXXXXXXXXXXXXXXX2
            : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX7, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX8 : out std_logic;  MXXXXXXXXXXXXXXXXXX3
            : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX10 : out std_logic;  
            MXXXXXXXXXXXXXXXXXX4 : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXXXX11
            : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXX1 : in std_logic;  
            MXXXXXXXXXXXXXXFXWXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXXXXX :
            in std_logic;  MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX : out 
            std_logic;  MXMXXXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXX3, XXXXXXXXXXXX 
            : in std_logic;  MXXXXXXXXXXXXXXXXXXPXXXXXXXX, XXXXXXX, XFXXXXXXXXX
            : out std_logic;  MXXXXXXXXXXXXXXYXXXX, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, MXMXXXXXXXXXXXXXXX3, XFXXXXXXXXXXX, 
            MXMXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXXXX5
            , MXXXXXXXXXXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX6, 
            MXXXXXXXXXXXXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXXXX7, 
            MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXMXMPXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXXXXXXMXMPXXXX, MXXXXXXXXXXXXXXXXXXXMXMPXXXX0, 
            MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXPXXXX : out std_logic;  MXMXXXXXXXXXXXXXXX10 : 
            in std_logic;  MXXXXXXXXXXXXXXXXXX6 : out std_logic;  XXMXXXXX : in
            std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0 : in 
            std_logic;  MXXXXXXXXXXXXXXXXXX7 : out std_logic;  XXXXXXXX : in 
            std_logic;  MXXXXXXXXXXXXXXXXXX8 : out std_logic;  XXXXXXXX0 : in 
            std_logic;  MXXXXXXXXXXXXXXXXXX9 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXXXXXX10, 
            MXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXX13
            : out std_logic;  MXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXX0 : 
            in std_logic;  XXMXXXX : out std_logic_vector (7 downto 0);  
            MXXXXXXXXXXXXXXYXXXX0, MXXXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXVXXXXXX, XXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXX2, 
            XXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1 : 
            in std_logic;  MXXXXXXXXXXXXXXXXXXXXXVXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXXVXX, MXXXXXXXXXXXXXXXXXXXXXXXVXX0, 
            MXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXX5 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXPXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXXXXX7, 
            MXXXXXXXXXXXXXXXXXXXXXXX8 : in std_logic;  MXXXXXXXXXXXXXXXXXX14 : 
            out std_logic;  MXXXXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXXXFXWXXX, 
            MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, MXXXXXXXXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXXXX11 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXFXXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXWXXX, MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0, 
            XXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXFXWXXX0
            : in std_logic;  XFXXXXXX : out std_logic_vector (8 downto 3);  
            MXXXXXXXXXXXXXPXHXXXXXX : in std_logic;  XXMXXXXX0 : out 
            std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXPXHXXXXXX0, 
            MXXXXXXXXXXXXXPXHXXXXXX1, MXXXXXXXXXXXXXPXHXXXXXX2, 
            MXXXXXXXXXXXXXPXHXXXXXX3, MXXXXXXXXXXXXXPXHXXXXXX4, 
            MXXXXXXXXXXXXXPXHXXXXXX5, MXXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXFXWXXX1, 
            MXXXXXXXXXXXXXPXHXXXXXX6, MXXXXXXXXXXXXXXXXXXFXWXXX2, 
            MXXXXXXXXXXXXXMXMPXXXXXXX1, MXXXXXXXXXXXXXXYXXXX1, 
            MXXXXXXXXXXXXXXXXXXX6, XXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX1 :
            in std_logic;  MXXXXXXXXXXXXXXXXXXX7 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  XFXXXXXXXXXXXXXXXXX, 
            XFXXXXXXXXXXXXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXMXMXMXXXX, 
            MXMXXXXXXXXXXXXXXX12, MXMXXXXXXXXXXXXXXX13, MXMXXXXXXXXXXXXXXX14, 
            MXMXXXXXXXXXXXXXXX15 : in std_logic;  MXXXXXXXXXXXXXXFXXXXXXXXX : 
            out std_logic;  MXXXXXXXXXXXXXXXMXXX, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX, MXXXXXXXXXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0
            , MXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX, 
            MXXXXXXXXXXXXXXXMXXX0, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2, MXXXXXXXXXXXXXXXXXXMXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3
            , MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXPXLXXXXXX, MXXXXXXXXXXXXXPXLXXXXXX0, 
            MXXXXXXXXXXXXXPXLXXXXXX1, MXXXXXXXXXXXXXPXLXXXXXX2, 
            MXXXXXXXXXXXXXPXLXXXXXX3, MXXXXXXXXXXXXXPXLXXXXXX4, 
            MXXXXXXXXXXXXXPXLXXXXXX5, MXXXXXXXXXXXXXXXXXX18, 
            MXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX0, MXXXXXXXXXXXXXXYXXXXXX, 
            MXXXXXXXXXXXXXXXXXXX10 : in std_logic;  XXMXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXX7, 
            MXMXXXXXXXXXXXXXXX16, MXMXXXXXXXXXXXXXXX17, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXX2, MXXXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXPXXXXXXX : in std_logic;  XFXXXXXX0 : in 
            std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXMXXX, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXPXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXPXXXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXPXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXX, MXXXXXXXXXXXXXXFXXXXXPXXXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXXX4, XFXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXMXXX1, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1, 
            MXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3, 
            MXXXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXFXXXXXXLXXXX2, 
            MXXXXXXXXXXXXXXXMXXX2, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2, 
            MXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXYXXXX2, MXXXXXXXXXXXXXXYXX, 
            MXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXMXMPXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXMXXX0, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8, MXXXXXXXXXXXXXPXLXXXXXX6, 
            MXXXXXXXXXXXXXXXXXX21, MXMXXXXXXXXXXXXXXX18, MXMXXXXXXXXXXXXXXX19 :
            in std_logic;  MXXXXXXXXXXXXXXXXXX22, XFXWX : out std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5, MXXXXXXXXXXXXXXFXXXXXXXXXXXX5,
            MXXXXXXXXXXXXXXFXXXXXXLXXXX3, MXXXXXXXXXXXXXXFXXXXXXXMXXX0, 
            MXXXXXXXXXXXXXXXXXX23, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7, MXXXXXXXXXXXXXXXMXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3, MXXXXXXXXXXXXXXXXXXMXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9, MXXXXXXXXXXXXXXXXXXXHXXX, 
            MXXXXXXXXXXXXXXXXXXFXWX, MXXXXXXXXXXXXXXXMXXX4, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4, MXXXXXXXXXXXXXXXXXXMXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11, MXXXXXXXXXXXXXXXXXXXHXXX0, 
            MXXXXXXXXXXXXXXXMXXX5, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2, MXXXXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXX3, MXMXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXX3,
            MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX4,
            MXXXXXXXXXXXXXXFXXXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12, MXXXXXXXXXXXXXXXXXX24, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12, MXXXXXXXXXXXXXXFXXXXXXLXXXX4,
            MXXXXXXXXXXXXXXXMXXX6, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXX4, MXMXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXX5,
            MXMXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXYXX0, MXXXXXXXXXXXXXXXXXX25, 
            MXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXX9 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXPXXXXXX0 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXX11, 
            MXXXXXXXXXXXXXXXXXX26, MXXXXXXXXXXXXXXXXXXXXX12, 
            MXXXXXXXXXXXXXXXXXXXXX13 : in std_logic;  XXMWX, XFXXX : out 
            std_logic;  MXXXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXXXX15 : in
            std_logic);
   end component;
   
   component XYXX0002
      port( MXXXXXXXXXXXXXXXXXXXFXWXXX, MXXXXXXXXXXXXXXXXXXFXWXXX : out 
            std_logic;  MXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, XLXXPX, MXXXXXXXXXXXXXXXXXXXXXXXX 
            : in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX : out std_logic;  ramaddr 
            : in std_logic_vector (5 downto 3);  XFXXXXXXXXXX, XFXXXXXXXXXXXX :
            in std_logic;  MXXXXXXXXXXXXXXXXXXFXWXXX0 : out std_logic;  
            MXXXXXXXXXXXXXXYXX, MXXXXXXXXXXXXXMXMPXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX, 
            MXXXXXXXXXXXXXMXMPXXXXXX : in std_logic;  MXMPXXXXWXXX : out 
            std_logic;  MXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXYXXXXXX, MXXXXXXXXXXXXXMXMPXXXXXXX0, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX0 : in 
            std_logic;  MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXFXWXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXX : in std_logic;  MXMPXXX : out std_logic;  
            XFXXXXXXXXXX0, XFXXXXXXXXXX1 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXFXWXXXXX : out std_logic;  XXXXXPXXX : in 
            std_logic;  MXXXXXXXXXXXXXXXMXMXXXLXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXYXXXX, MXXXXXXXXXXXXXXXXXXXXXXXVXX, 
            MXXXXXXXXXXXXXXXXXFXXXHX, MXXXXXXXXXXXXXXXXXXLLXX, 
            MXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX0, 
            MXXXXXXXXXXXXXPXLXXXXXX1 : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX1 
            : in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX2 : out std_logic;  
            XXXXXXXX : in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX3 : out std_logic;
            MXXXXXXXXXXXXXXXXXXXXX2 : in std_logic;  MXXXXXXXXXXXXXPXLXXXXXX4 :
            out std_logic;  XXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXX3 : in std_logic; 
            MXXXXXXXXXXXXXPXHXXXXXX, MXXXXXXXXXXXXXPXHXXXXXX0 : out std_logic; 
            MXMXXXX : out std_logic_vector (15 downto 0);  XXXXXXXX1, XXXXXXXX2
            , MXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXXXVXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXVXXXXXX2, MXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXVXXXXXX3, MXXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXPXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXX4, MXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXHXXX, MXXXXXXXXXXXXXXXXXXXHXXX0, 
            MXXXXXXXXXXXXXXXXXXXHXXX1, MXXXXXXXXXXXXXXXXXXXXX4, 
            MXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX6, XXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXX7, MXMXXXX0, MXXXXXXXXXXXXXXXXXXX8, 
            MXXXXXXXXXXXXXXXXVXLXX, MXXXXXXXXXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXYXXXX0, 
            MXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXX12, 
            MXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXXXXXX2 : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0
            , MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2, MXXXXXXXXXXXXXXXXXXFXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11, 
            MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12 : out std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXWXXX, 
            MXXXXXXXXXXXXXXFXWXXX : in std_logic;  XXMXXXXX : in 
            std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXXFXXXXXMXXXXX : out 
            std_logic;  MXMXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXX0 : in std_logic;
            MXXXXXXXXXXXXXPXHXXXXXX1, MXXXXXXXXXXXXXPXHXXXXXX2, 
            MXXXXXXXXXXXXXPXHXXXXXX3, MXXXXXXXXXXXXXPXHXXXXXX4, 
            MXXXXXXXXXXXXXPXLXXXXXX5 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXFXWXXX1, MXMXXXXXXXXXXXXXXX1, 
            MXMXXXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXXXX3 : in std_logic;  
            MXXXXXXXXXXXXXPXHXXXXXX5, MXXXXXXXXXXXXXPXHXXXXXX6, 
            MXXXXXXXXXXXXXPXLXXXXXX6 : out std_logic;  MXXXXXXXXXXXXXXYXX0, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXX0, MXXXXXXXXXXXXXMXMPXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXJXMP, 
            MXXXXXXXXXXXXXXXXXXX15 : in std_logic;  MXXXXXXXXXXXXXXXXXMXVXWXXX 
            : out std_logic;  MXXXXXXXXXXXXXXXXXXX16, 
            MXXXXXXXXXXXXXMXMPXXXXXXX2, MXXXXXXXXXXXXXXXXXXXX0 : in std_logic; 
            MXXXXXXXXXXXXXXXXXXFXWXXX2 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXWXXX0, MXMXXXXXXXXXXXXXXX4, 
            MXMXXXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXFXXXHX
            : in std_logic;  MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX : out 
            std_logic;  MXXXXXXXXXXXXXXYXXXX1, MXXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX, 
            MXXXXXXXXXXXXXXXXXXLL : in std_logic;  MXMXXXXX : in 
            std_logic_vector (7 downto 0);  MXMXXXXXXXXXXXXXXX7, 
            MXXXXXXXXXXXXXXXXXXXPXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, 
            XFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXXXXX, MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX9
            , MXMXXXXXXXXXXXXXXX10, MXMXXXXXXXXXXXXXXX11, MXMXXXXXXXXXXXXXXX12,
            MXMXXXXXXXXXXXXXXX13, MXMXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXX18,
            MXXXXXXXXXXXXXXYFLXX, MXXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXYXX1 :
            in std_logic;  MXXXXXXXXXXXXXXXXXXPXXLXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX4, XXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX2, 
            MXMXXXXXXXXXXXXXXX15, MXMXXXXXXXXXXXXXXX16, MXMXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX5 : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXFXWXXX0 : out std_logic;  XFXWX, 
            MXXXXXXXXXXXXXXXXXX : in std_logic;  MXXXXXXXXXXXXXXXXXXMXMPXXXX : 
            out std_logic;  MXXXXXXXXXXXXXXXXXXX21, XXMXXXXXXX, 
            MXXXXXXXXXXXXXMXMPXXXXX, XXXXXXXX3, MXXXXXXXXXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXXXXFXXXHXXX, MXXXXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXX0
            , MXXXXXXXXXXXXXXFXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXX6 : in std_logic;  
            MXXXXXXXXXXXXXXXMXMXMXXXX, MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, 
            MXMWXXXXXX, MXXXXXXXXXXXXXMXMXXXX, MXMXX : out std_logic;  XFXXXXXX
            : in std_logic_vector (7 downto 0);  MXXXXXXXXXXXXXXXXXXXXX7, 
            MXMXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXX3, 
            MXMXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXX6, 
            MXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXX11, 
            MXXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXXX13, 
            MXXXXXXXXXXXXXXXXXXXXX14 : in std_logic);
   end component;
   
   component XYXX0001
      port( MXXXXXXXXXXXXXMXMXXXX, XLXXPX, MXXXXXXXXXXXXXXXXXXXXXX : in 
            std_logic;  MXXXXXXXXXXXXXXXXXXXXX, XXXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXX0 : in std_logic;  XXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXXXX0, XXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXX1, 
            XXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXX2 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX, MXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXWXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXXXXXXXWXXX : out std_logic;  MXXXXXXXXXXXXXXYXX, 
            MXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXX3
            , MXXXXXXXXXXXXXXXXXXFXWXXXXX, XFXXXXXXXXXX, XFXXXXXXXXXX0, 
            MXXXXXXXXXXXXXMXMPXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXVXX, 
            MXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXX7
            , MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX8, XFXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXX10, 
            MXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXX12, 
            MXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXMXMPXXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXXXX6, 
            MXXXXXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, 
            MXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXX17, 
            MXXXXXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXXXXXX19, 
            MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXXXX7, 
            MXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXX20, 
            MXXXXXXXXXXXXXXXXXXXXXXVXX0, MXXXXXXXXXXXXXXYXXXX, 
            MXXXXXXXXXXXXXXXXXXX21 : in std_logic;  
            MXXXXXXXXXXXXXXXXXPXWXXXXWXXX : out std_logic;  XFXXXXXXXXXX1, 
            MXXXXXXXXXXXXXXXXXXFXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXX, 
            MXXXXXXXXXXXXXXYXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0
            , MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXFXWXXX, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXX, MXXXXXXXXXXXXXXXXXXX23, 
            MXXXXXXXXXXXXXXXXXXPXXXXXXXX, MXXXXXXXXXXXXXXYXXXX1, 
            MXXXXXXXXXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXXXX25, 
            MXXXXXXXXXXXXXXXXXXX26, MXXXXXXXXXXXXXXXXXXX27, 
            MXXXXXXXXXXXXXXXXXXX28, MXXXXXXXXXXXXXXXXXXXXX9, 
            MXXXXXXXXXXXXXXXXXXX29 : in std_logic;  MXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXX8, 
            MXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXX10 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXX30, MXXXXXXXXXXXXXXXXXXXXXXXVXX0, 
            MXXXXXXXXXXXXXXXXXX11, MXMXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXX12, 
            MXXXXXXXXXXXXXXXXXX13 : in std_logic;  MXXXXXXXXXXXXXXXXXX14 : out 
            std_logic;  MXMXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX1, 
            MXMXXXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXXXX3, MXMXXXXXXXXXXXXXXX4, 
            MXMXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXXYXXXX2,
            MXXXXXXXXXXXXXMXMPXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXXXXXX32, MXXXXXXX : in std_logic;  
            MXXXXXXXXXXXXXXXXLXXXXXXX, MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX,
            MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXX11, 
            MXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXVXX, 
            MXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXX33, 
            MXXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXXXX : in 
            std_logic;  MXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXX0, 
            MXXXXXXXXXXXXXXYFLXX : out std_logic;  MXXXXXXXXXXXXXXXXXXXXX12 : 
            in std_logic;  MXMXXXXX : out std_logic_vector (7 downto 0);  
            MXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, 
            MXXXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXFXXXXXXXXXX0 : in 
            std_logic;  MXXXXXXXXXXXXXXXMXXX : out std_logic;  
            MXXXXXXXXXXXXXXFXXXXXXXXXX1 : in std_logic;  MXXXXXXXXXXXXXXXMXXX0,
            MXXXXXXXXXXXXXXXMXXX1, MXXXXXXXXXXXXXXXMXXX2 : out std_logic;  
            MXMXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, 
            MXMXXXXXXXXXXXXXXX7, MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX9, 
            MXMXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXX34, 
            MXXXXXXXXXXXXXXXXXXX35, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, 
            MXXXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXXX4, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2, MXXXXXXXXXXXXXXXXXXXXXXXVXX1, 
            MXXXXXXXXXXXXXXXXXXXXX15 : in std_logic;  
            MXXXXXXXXXXXXXXXXLXXXXXXX0 : out std_logic;  MXXXXXXXXXXXXXXXXXXX36
            , MXXXXXXXXXXXXXXXXXXX37, MXMXXXXXXXXXXXXXXX11, 
            MXXXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXXXXXXVXX2, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, MXXXXXXXXXXXXXXXXXXX38, 
            MXXXXXXXXXXXXXXXXXXX39, MXXXXXXXXXXXXXXXXXXX40, 
            MXXXXXXXXXXXXXXXXXXXXXXXVXX3, MXXXXXXXXXXXXXXXXXXXX5, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX2 : in std_logic;  MXXXXXXXXXXXXXXXMXXX3 
            : out std_logic;  XFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX3, 
            MXXXXXXXXXXXXXXFXXXXXXXXXX4 : in std_logic;  ramaddr : in 
            std_logic_vector (6 downto 1);  MXXXXXXXXXXXXXXXMXXX4, 
            MXXXXXXXXXXXXXXXMXXX5 : out std_logic;  MXXXXXXXXXXXXXXYXXXXXX, 
            MXXXXXXXXXXXXXMXMPXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXX2, 
            MXXXXXXXXXXXXXXYXX0 : in std_logic;  MXXXXXXXXXXXXXXXXXVXXXXXX, 
            MXXXXXXXXXXXXXXXXXXXXXXWXXX0, MXXXXXXXXXXXXXXXXXXXXXXWXXX1, 
            MXXXXXXXXXXXXXXXMXXX6, MXXXXXXXXXXXXXXXJXMP, MXXXXXXXXXXXXXXXXVXLXX
            : out std_logic;  MXXXXXXXXXXXXXXXXXXXX6, MXMXXXXXXXXXXXXX0, 
            MXMXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX7, 
            MXXXXXXXXXXXXXXFXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXX8, 
            MXXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXXX10 : in std_logic;  
            MXXXXXXXXXXXXXXXXLXXXXXXX1 : out std_logic;  
            MXXXXXXXXXXXXXXXXXXXX11 : in std_logic;  MXXXXXXXXXXXXXXXXLXXXXXXX2
            : out std_logic;  MXXXXXXXXXXXXXXXXXXXX12, 
            MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX : in std_logic);
   end component;
   
   signal port0o0_7_port, port0o0_6_port, port0o0_5_port, port0o0_4_port, 
      port0o0_3_port, port0o0_2_port, port0o0_1_port, port0o0_0_port, 
      port1o0_7_port, port1o0_6_port, port1o0_5_port, port1o0_4_port, 
      port1o0_3_port, port1o0_2_port, port1o0_1_port, port1o0_0_port, 
      port2o0_7_port, port2o0_6_port, port2o0_5_port, port2o0_4_port, 
      port2o0_3_port, port2o0_2_port, port2o0_1_port, port2o0_0_port, 
      port3o0_7_port, port3o0_6_port, port3o0_5_port, port3o0_4_port, 
      port3o0_3_port, port3o0_2_port, port3o0_1_port, port3o0_0_port, 
      memdatao0_7_port, memdatao0_6_port, memdatao0_5_port, memdatao0_4_port, 
      memdatao0_3_port, memdatao0_2_port, memdatao0_1_port, memdatao0_0_port, 
      memaddr0_15_port, memaddr0_14_port, memaddr0_13_port, memaddr0_12_port, 
      memaddr0_11_port, memaddr0_10_port, memaddr0_9_port, memaddr0_8_port, 
      memaddr0_7_port, memaddr0_6_port, memaddr0_5_port, memaddr0_4_port, 
      memaddr0_3_port, memaddr0_2_port, memaddr0_1_port, memaddr0_0_port, 
      ramaddr0_7_port, ramaddr_6, ramaddr_5, ramaddr_4, ramaddr_3, ramaddr_2, 
      ramaddr_1, ramaddr_0, sfrdatao0_7_port, sfrdatao0_6_port, 
      sfrdatao0_5_port, sfrdatao0_4_port, sfrdatao0_3_port, sfrdatao0_2_port, 
      sfrdatao0_1_port, sfrdatao0_0_port, nrsto0, nrsto_nc0, clkcpu_en0, 
      clkper_en0, sfrwe0, TrigOut0, XXXXXX8, XXXXXX9, XXXXXXXXXX6, XXXXXXXXXX7,
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, XXXXXXXXX1, 
      MXMXXXXXXXXXXXXXXXXX, XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, 
      MXMXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXXXX2, XXXXXXXXXXXXXXXXXX, XXXXXXXXXX8, XXXXXXXXXX9, 
      XXXXXXXXX2, XXXXXX10, MXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXLXXXXXXX, MXXXXXXX4, MXMPXXXXWXXX, XXXXXXXXXX10, 
      XXXXXX11, XXXXXXXXXX11, MXXXXX6, MXXXXXXXXXXXXXXXXLXXXXXXX0, 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1, MXMXXXXXXXXXXXXXXX, 
      XXXXXXXX11, MXXXXXX1, XXXXXX12, XXX10, XXXXXX13, XXXXXX14, XXXXXX15, 
      XXXXXXX24, MXXX16, XXXXXX16, MXXXXX7, XXXXXXXXX3, 
      MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, 
      MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX, MXXXXXXX5, XXX11, XXXX17, XXXX18,
      XXXXXXXX12, XXXXXXXX13, XXXXXXXXXX12, XXXXXXXXXXXXXX, XXXXXXXXXXXX3, 
      XXXXXXXX14, XXXXXXXXX4, MXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXX1, 
      MXXXXX8, MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2, MXMXXXXXXXXXXXXX, MXXXXXX2, 
      XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3, MXMXXXXXXXXXXXXX0, 
      XXXXXXXXXX13, MXXXXX9, MXXXXXXXXXXXXXXXPMXXXXXXXXLXXX, XXXXX31, XXXXX32, 
      XFXXXXXXXXXX, XFXXXXXXXXXXXX, XXXXX33, XXXXX34, XXXXX35, MXXXXX10, 
      XXXXXXX25, MXXXXX11, XXXX19, XXXXXX17, 
      MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, XXXXXXX26, MXXX17, MXXXX12, 
      XXXXXXX27, MXXXX13, MXXXXX12, MXXXXXXXXXXXXXXXXXFXXXHXXX, XXXXXXXX15, 
      XXXXXXXX16, XXXXXXXX17, MXXXX14, XXXXX36, XFXXXXXXXXXXX, XFXXXXXXXXXXX0, 
      MXMXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXXXX2, 
      MXMXXXXXXXXXXXXXXX3, MXMXXXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXXXX5, 
      MXMXXXXXXXXXXXXXXX6, XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4, 
      MXMXXXXXXXXXXXXXXX7, MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX9, 
      MXMXXXXXXXXXXXXXXX10, MXMXXXXXXXXXXXXXXX11, MXMXXXXXXXXXXXXXXX12, 
      MXMXXXXXXXXXXXXXXX13, MXMXXXXXXXXXXXXXXX14, MXXXXX13, MXXXXX14, 
      XXXXXXXX18, MXMXXXXXXXXXXXXXXX15, MXMXXXXXXXXXXXXXXX16, 
      MXMXXXXXXXXXXXXXXX17, XXXXXXX28, XXXXXXXXXX14, XXXXXXX29, 
      MXMXXXXXXXXXXXXXXX18, MXMXXXXXXXXXXXXXXX19, MXMXXXXXXXXXXXXXXX20, 
      XXXXXXXXXXXXXXXX0, XXXXXXXXXX15, MXXXXXXXXXXXXXXXXXFXXXHX, 
      MXXXXXXXXXXXXXXXXXXFXXXHX, XXXXXXMXXX, XXXXXXXXXX16, MXXXXX15, 
      MXXXXXXXXXXXXXMXMPXXXXXX, MXXXXXX3, MXXXXXXX6, XXXXXPXXX, MXXXXX16, 
      MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX, 
      MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXXXX1, 
      MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, 
      MXXXXX17, MXXXXX18, MXXXXX19, MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXX, 
      XFXXXXXXXXXX0, XFXXXXXXXXXX1, XXXXXXXXXX17, XXXXXXX30, XXXXXXXX19, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX36, MXXX18, XXXXXXXXXXXX4, 
      XXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXLXXXXXXX2, 
      MXXXXXXXX, MXXXXXX4, MXXXXXX5, MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX, 
      MXXXXXXX7, MXXXXX20, XXXXXXXXXX18, XXXXXXX31, MXXXXXXXXXXXXXXXXXXX0, 
      MXXXXXXX8, MXXXXXX6, MXXXXXXX9, MXXX19, MXXXXX21, MXXXXX22, XXXXXX18, 
      MXXXXX23, MXX5, XXXXXXXXX5, MXXXXXXX10, MXXXX15, MXXXXXXX11, MXXXXX24, 
      MXXXXXXX12, XXXXXXXX20, XXXXXXX32, MXXXXX25, XXXXXXXXXXXX5, XXXXXXX33, 
      MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX, XFXXXXXXXXXXXXXXXXX, XXXXXXXXXXXX6, 
      MXXXXXXXXXXXXXXXXXXXXXXX4, XXXXXXXX21, XFXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXXXXXXXX5, XFXXXXXXXXXXXXXXXXX0, MXXXXX26, XXXXXXX34, 
      XXXXXXXXX6, MXXXXX27, MXXXXX28, MXXXXXX7, MXXXXXXX13, MXXXXXXXX0, 
      MXXXXXX8, MXXXXXX9, MXXXXX29, MXXXXXXX14, XXXXXXXXX7, MXXXXXX10, 
      MXMXXXXXXXXXXXXX1, XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5, MXXXXX30, 
      XXXXXXXXXX19, XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6, 
      MXMXXXXXXXXXXXXX2, XXXXXXX35, XXXXXXXXXX20, XXX12, MXXX20, 
      MXXXXXXXXXXXXXXXXXFXXXHX0, MXMXXXXXXXXXXXXX3, MXMXXXXXXXXXXXXX4, 
      MXMXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXX6, JXXXXX, XXXXXXXXXXX, MXMWXXXXXX0, 
      XXXXXPXWX, XXXXXXXX22, XXXXXXXX23, XXXXXXXX24, XXXXXXXX25, 
      MXXXXXXXXXXXXXXXXXXXXXXX6, XXXXXXXXP, XXXXXXXX26, XXXXXXXX27, URSTB, 
      UDRCK, UDRCK_1, XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX1, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX2, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX3, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX4, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX5, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX6, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXP, 
      XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXPX, 
      MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXX7, 
      MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXX8, 
      MXXXXXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2,
      MXXXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXPXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX, MXXXXXXXXXXXXXXXPXXXXXXXXX, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX0, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX1, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX2, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX3, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX4, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX5, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX6, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX7, 
      MXXXXXXXXXXXXXXXPXXXXXXXXX0, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX8, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX9, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX10, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX11, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX12,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX13, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX14,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX15, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX16,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX17, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX18,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX19, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX20,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX21, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX22,
      MXXXXXXXXXXXXXXXPXXXXXXXXXX0, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX23, 
      MXXXXXXXXXXXXXXXPXXXXXXXXXX1, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX24, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX25, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX26,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX27, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX28,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX29, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX30,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX31, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX32,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX33, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX34,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX35, MXXXXXXXXXXXXXXXPXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, MXXXXXXXXXXXXXXXPXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXPXXXXXXXXX2, MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX3, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX5, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX6, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX7, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX8, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX9, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX10, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX11, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX12, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX13, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX14, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX15, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX16, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX17, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX18, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX19, 
      MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, 
      MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX20, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX21, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX36, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX37,
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX38, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX22, 
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX23, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX39, MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX40,
      MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX24, 
      MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX41, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX3, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX5, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXX, MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXFF, MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXPMXXXXXXX, 
      MXXXXXXXXXXXXXXXPMXXXXXXX0, MXXXXXXXXXXXXXXXPMXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXPMXXXXXXXXXXX2, MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXX, 
      MXXXXXXXXXXXXXXXPMXXXXXXXLXXPXXXXXXXPXXXX, 
      MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXXXPXXXX, 
      MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXXXPXXXX, 
      MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, 
      MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX, MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX0
      , MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX1, MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX
      , MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX0, MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX1, MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX3, 
      MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX2, MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX5, MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX3, 
      MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXLXXXXLXXXMXXXXXXX, MXXXXXXXXXXXXXXXXLXXXXLXXXMXXXXXXX0, 
      MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX6, MXXXXXXXXXXXXXXXXLXXXXLXXXXX, 
      MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX4, XXXXXXXXXXXXXXXXXJXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX37, 
      MXXXXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXX13, 
      MXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, 
      MXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX38, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX15, MXXXXXXXXXXXXXXXXXXX7, 
      MXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXXX7, 
      MXXXXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXXXX9, 
      MXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXX9
      , MXXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXX10, 
      MXXXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXXXX14, 
      MXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXLXXXXXXXXXX, 
      MXXXXXXXXXXXXXXLXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, 
      MXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXX15, 
      MXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXX17, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXX, MXXXXXXXXXXXXXXXXXXX18, 
      MXXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXX20, 
      MXXXXXXXXXXXXXXXXXXX21, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX18, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXX16, 
      MXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXX23,
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX6, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX7, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXXX24, 
      MXXXXXXXXXXXXXXXXXXX25, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX19, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXXXX26, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX39, MXXXXXXXXXXXXXXXXXXX27, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXX28, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXX29, 
      MXXXXXXXXXXXXXXXXXXX30, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX11, 
      MXXXXXXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXXXXXXX32, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX21, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX12, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX13, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXX33, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXX34, 
      MXXXXXXXXXXXXXXXXXXX35, MXXXXXXXXXXXXXXXXXXX36, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX23, MXXXXXXXXXXXXXXXXXXX37, 
      MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX38, 
      MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1,
      MXXXXXXXXXXXXXXXXXXX39, MXXXXXXXXXXXXXXXXXXX40, MXXXXXXXXXXXXXXXXXXX41, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX24, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX15, MXXXXXXXXXXXXXXXXXXXXXXX14, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX25, MXXXXXXXXXXXXXXXXXXPXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXX42, 
      MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX5, 
      MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXX43, 
      MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXX44, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX26, MXXXXXXXXXXXXXXXXXXX45, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXX46, 
      MXXXXXXXXXXXXXXXXXXX47, MXXXXXXXXXXXXXXXXXXX48, MXXXXXXXXXXXXXXXXXXX49, 
      MXXXXXXXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXXXXXX50, MXXXXXXXXXXXXXXXXXXX51,
      MXXXXXXXXXXXXXXXXXXXXXXVXX, MXXXXXXXXXXXXXXXXXXX52, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXXXXXXXXXXVXX0, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXXXXXXVXX2, 
      MXXXXXXXXXXXXXXXXXXX53, MXXXXXXXXXXXXXXXXXXX54, MXXXXXXXXXXXXXXXXXXX55, 
      MXXXXXXXXXXXXXXXXXXXXXXVXX0, MXXXXXXXXXXXXXXXXXXX56, 
      MXXXXXXXXXXXXXXXXXXX57, MXXXXXXXXXXXXXXXXXXXXXXXVXX3, 
      MXXXXXXXXXXXXXXXXXXX58, MXXXXXXXXXXXXXXXXXXX59, MXXXXXXXXXXXXXXXXXXX60, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXX4, MXXXXXXXXXXXXXXXXXXX61, 
      MXXXXXXXXXXXXXXXXXXX62, MXXXXXXXXXXXXXXXXXXX63, MXXXXXXXXXXXXXXXXXXX64, 
      MXXXXXXXXXXXXXXXXXXX65, MXXXXXXXXXXXXXXXXXXPXXXXXXXX, 
      MXXXXXXXXXXXXXXLXXXXXXXXXX0, MXXXXXXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXX15, 
      MXXXXXXXXXXXXXXXXXXX66, MXXXXXXXXXXXXXXXXXXX67, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXMXXX, MXXXXXXXXXXXXXXXXXXXXX19, 
      MXXXXXXXXXXXXXXXXXXX68, MXXXXXXXXXXXXXXXXXXX69, MXXXXXXXXXXXXXXXXXXXXX20,
      MXXXXXXXXXXXXXXLXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXLXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXX70, MXXXXXXXXXXXXXXXXXXX71, MXXXXXXXXXXXXXXXXXXXXX21,
      MXXXXXXXXXXXXXXXXXXPXXXXXX0, MXXXXXXXXXXXXXXXXXXX72, 
      MXXXXXXXXXXXXXXXXXXX73, MXXXXXXXXXXXXXXXXXXXXXXX16, 
      MXXXXXXXXXXXXXXXXXXX74, MXXXXXXXXXXXXXXXXXXX75, MXXXXXXXXXXXXXXXXXXX76, 
      MXXXXXXXXXXXXXXXXXXX77, MXXXXXXXXXXXXXXXXXXX78, MXXXXXXXXXXXXXXXXXXX79, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, MXXXXXXXXXXXXXXXXXXX80, 
      MXXXXXXXXXXXXXXXXXXX81, MXXXXXXXXXXXXXXXXXXX82, MXXXXXXXXXXXXXXXXXXX83, 
      MXXXXXXXXXXXXXXXXXXX84, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2, 
      MXXXXXXXXXXXXXXXXXXX85, MXXXXXXXXXXXXXXXXXXX86, MXXXXXXXXXXXXXXXXXXX87, 
      MXXXXXXXXXXXXXXXXXXX88, MXXXXXXXXXXXXXXXXXXX89, MXXXXXXXXXXXXXXXXXXX90, 
      MXXXXXXXXXXXXXXXXXXX91, MXXXXXXXXXXXXXXXXXXX92, MXXXXXXXXXXXXXXXXXXX93, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXX3, 
      MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXX94, MXXXXXXXXXXXXXXXXXXX95,
      MXXXXXXXXXXXXXXXXXXX96, MXXXXXXXXXXXXXXXXXXX97, MXXXXXXXXXXXXXXXXXXX98, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXX5, MXXXXXXXXXXXXXXXXXXXXXXXVXX6, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXXVXX7, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXX8, MXXXXXXXXXXXXXXXXXXXXXXXVXX9, 
      MXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXX99, 
      MXXXXXXXXXXXXXXXXXXX100, MXXXXXXXXXXXXXXXXXXXXX23, 
      MXXXXXXXXXXXXXXXXXXX101, MXXXXXXXXXXXXXXXXXXX102, 
      MXXXXXXXXXXXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXXXX103, 
      MXXXXXXXXXXXXXXXXXXX104, MXXXXXXXXXXXXXXXXXXX105, MXXXXXXXXXXXXXXXXXXX106
      , MXXXXXXXXXXXXXXXXXXX107, MXXXXXXXXXXXXXXXXXXX108, 
      MXXXXXXXXXXXXXXXXXXX109, MXXXXXXXXXXXXXXXXXXX110, MXXXXXXXXXXXXXXXXXXX111
      , MXXXXXXXXXXXXXXXXXXX112, MXXXXXXXXXXXXXXXXXXXXXXXVXX10, 
      MXXXXXXXXXXXXXXXXXXX113, MXXXXXXXXXXXXXXXXXXXXXXXVXX11, 
      MXXXXXXXXXXXXXXXXXXX114, MXXXXXXXXXXXXXXXXXXXXX25, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXX4, MXXXXXXXXXXXXXXXXXXX115, 
      MXXXXXXXXXXXXXXXXXXXXX26, MXXXXXXXXXXXXXXXXXXXXX27, 
      MXXXXXXXXXXXXXXXXXXX116, MXXXXXXXXXXXXXXXXXXX117, 
      MXXXXXXXXXXXXXXXXXXXXXXXVXXXX5, MXXXXXXXXXXXXXXXXXXX118, 
      MXXXXXXXXXXXXXXXXXXX119, MXXXXXXXXXXXXXXXXXXXXXXXVXXXX6, 
      MXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXLXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXLXXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXLXXXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXXXXXX28, MXXXXXXXXXXXXXXLXXXXXXXXXXXX3, 
      MXXXXXXXXXXXXXXXXXXX120, MXXXXXXXXXXXXXXXXXXX121, 
      MXXXXXXXXXXXXXXXXXXXXXVXX, MXXXXXXXXXXXXXXXXXXX122, 
      MXXXXXXXXXXXXXXXXXXX123, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX27, 
      MXXXXXXXXXXXXXXXXXXXXX29, MXXXXXXXXXXXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXXX30, MXXXXXXXXXXXXXXXXXXXXXX0, 
      MXXXXXXXXXXXXXXLXXXVXX, MXXXXXXXXXXXXXXLXXXVX, 
      MXXXXXXXXXXXXXXXXXXXXXXXXLXX, MXXXXXXXXXXXXXXLXXXVX0, MXXXXXXXXXXXXXXXX1,
      MXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXFXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXX2, 
      MXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXX5, 
      MXXXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXXXX8, 
      MXXXXXXXXXXXXXXXXVXLXX, MXXXXXXXXXXXXXXXJXMP, MXXXXXXXXXXXXXXXXXXXXXXWXXX
      , MXXXXXXXXXXXXXXXXXXXXXXWXXX0, MXXXXXXXXXXXXXXYXX, 
      MXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXVXXXXXX, 
      MXXXXXXXXXXXXXMXMPXXXXXXX, MXXXXXXXXXXXXXXYXXXXXX, MXXXXXXXXXXXXXXXXXXXX9
      , MXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXYFLXX,
      MXXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXMXMPXXXXXXX0, MXXXXXXXXXXXXXXYXXXX
      , MXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXX7, 
      MXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXX10, 
      MXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXYXXXX0, MXXXXXXXXXXXXXXXXXXXFXWXXX,
      MXXXXXXXXXXXXXXYXXXX1, MXXXXXXXXXXXXXXXXXXFXXXXXXX, 
      MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, MXXXXXXXXXXXXXXYXXXX2, 
      MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXMXMPXXXXXXX1, 
      MXXXXXXXXXXXXXMXMPXXXXXXX2, MXXXXXXXXXXXXXXXXXXFXWXXXXX, 
      MXXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXYXX0, 
      MXXXXXXXXXXXXXXXXXXXXXXWXXX1, MXXXXXXXXXXXXXXFXWXXX, 
      MXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXX14, 
      MXXXXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXX17, 
      MXXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXXX15, 
      MXXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXMXMXXXX
      , MXXXXXXXXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXXXXXXXXX32, 
      MXXXXXXXXXXXXXXXXXXXXX33, MXXXXXXXXXXXXXXXXXXXXX34, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1, 
      MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3, 
      MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4, MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5, 
      MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6, MXXXXXXXXXXXXXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXMXXX, MXXXXXXXXXXXXXXXMXXX0, 
      MXXXXXXXXXXXXXXXMXXX1, MXXXXXXXXXXXXXXXMXXX2, MXXXXXXXXXXXXXXXMXXX3, 
      MXXXXXXXXXXXXXXXMXXX4, MXXXXXXXXXXXXXXXMXXX5, MXXXXXXXXXXXXXXXMXXX6, 
      MXXXXXXXXXXXXXXFXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXXXX35, 
      MXXXXXXXXXXXXXXXXXXXLX, MXXXXXXXXXXXXXMXMPXXXXX, 
      MXXXXXXXXXXXXXXXXXXFXWXXX, MXXXXXXXXXXXXXXMXX, MXXXXXXXXXXXXXXXXXX18, 
      MXXXXXXXXXXXXXXXXXXFXWX, MXXXXXXXXXXXXXXXXXXFXWXXX0, 
      MXXXXXXXXXXXXXXXXXXFXWXXX1, MXXXXXXXXXXXXXXXXXXFXXXXX, 
      MXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXFXXXXXXXXXX5, 
      MXXXXXXXXXXXXXXFXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXXXXXX7, 
      MXXXXXXXXXXXXXXFXXXXXXLXXXX, MXXXXXXXXXXXXXXFXXXXXXLXXXX0, 
      MXXXXXXXXXXXXXXFXXXXXXLXXXX1, MXXXXXXXXXXXXXXFXXXXXXLXXXX2, 
      MXXXXXXXXXXXXXXFXXXXXXLXXXX3, MXXXXXXXXXXXXXXFXXXXXXLXXXX4, 
      MXXXXXXXXXXXXXXXXXXXHXXX, MXXXXXXXXXXXXXXXXXXXHXXX0, 
      MXXXXXXXXXXXXXXXXXXXHXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXXX7, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXX8, MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXX10, MXXXXXXXXXXXXXXFXXXXXXXXXXX11, 
      MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXYXLXXXXXX, 
      MXXXXXXXXXXXXXXYXLXXXXXX0, MXXXXXXXXXXXXXXYXLXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXX36, MXXXXXXXXXXXXXXXXXXXXX37, 
      MXXXXXXXXXXXXXXMWXXXXX, MXXXXXXXXXXXXXXXXXXX124, MXXXXXXXXXXXXXXXXXXX125,
      MXXXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXXX21, MXXXXXXXXXXXXXXXXXXXXXPFF, 
      MXXXXXXXXXXXXXXXXXXLL, MXXXXXXXXXXXXXXXXXMXVXWXXX, 
      MXXXXXXXXXXXXXXXXXXPXXLXX, MXXXXXXXXXXXXXXYXX1, 
      MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXPXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXPXXXXXX0, 
      MXXXXXXXXXXXXXXXXXXXMXMPXXXX, MXXXXXXXXXXXXXXXXXXXMXMPXXXX0, 
      MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXX126
      , MXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXLLXX, 
      MXXXXXXXXXXXXXXMWXXXXXXX, MXXXXXXXXXXXXXXXXXXXX18, 
      MXXXXXXXXXXXXXXMWXXXXXXX0, MXXXXXXXXXXXXXXXXXXMXMPXXXX, 
      MXXXXXXXXXXXXXXXXPPMX, MXXXXXXXXXXXXXXXXXXXXXXX18, 
      MXXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXPXXXXXX1, 
      MXXXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXX19, 
      MXXXXXXXXXXXXXXYXLXXXX, MXXXXXXXXXXXXXXYXLXXXX0, MXXXXXXXXXXXXXXYXLXXXX1,
      MXXXXXXXXXXXXXXYXLXXXX2, MXXXXXXXXXXXXXXXXYXLXXXXX, 
      MXXXXXXXXXXXXXXXXYXLXXXXX0, MXXXXXXXXXXXXXXXXYXLXXXXX1, 
      MXXXXXXXXXXXXXXXXYXLXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXX8, 
      MXXXXXXXXXXXXXXFXXXXXXXXXX9, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1,
      MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3,
      MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5,
      MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7,
      MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9,
      MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10, MXXXXXXXXXXXXXXXXXXXXX38, 
      MXXXXXXXXXXXXXXXXXXXXX39, MXXXXXXXXXXXXXXXXXXXXX40, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXX41, 
      MXXXXXXXXXXXXXXXXXXXXX42, MXXXXXXXXXXXXXXXXXXXXX43, 
      MXXXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXXXXX21
      , MXXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXXX44, 
      MXXXXXXXXXXXXXXXXXX23, MXXXXXXXXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXXXX127, 
      MXXXXXXXXXXXXXXXXXX25, MXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXX4, 
      MXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXX26, MXXXXXXXXXXXXXXFX, 
      MXXXXXXXXXXXXXXXL, MXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXX27, 
      MXXXXXXXXXXXXXXFX0, MXXXXXXXXXXXXXXXXXXFXWXXX2, MXXXXXXXXXXXXXXXXXXXX23, 
      MXXXXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12, MXXXXXXXXXXXXXXXXPXXXXXXXX, 
      MXXXXXXXXXXXXXXXXPXXXXXXXX0, MXXXXXXXXXXXXXXXXVXXXXXX, 
      MXXXXXXXXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXXXVXXXXXX1, 
      MXXXXXXXXXXXXXXXXVXXXXXX2, MXXXXXXXXXXXXXXXXVXXXXXX3, 
      MXXXXXXXXXXXXXXXXPXXXXXXXX1, MXXXXXXXXXXXXXXXXPXXXXXXXX2, 
      MXXXXXXXXXXXXXXFXXXXXMXXXXX, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1, 
      MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3, 
      MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5, 
      MXXXXXXXXXXXXXXXXXXXXX45, MXXXXXXXXXXXXXXXXXXXXX46, 
      MXXXXXXXXXXXXXXXXXXXXX47, MXXXXXXXXXXXXXXXXXXXXX48, 
      MXXXXXXXXXXXXXXXXXXXXX49, MXXXXXXXXXXXXXXXXXXXXX50, 
      MXXXXXXXXXXXXXXXXXXXXX51, MXXXXXXXXXXXXXXXXXXXXX52, 
      MXXXXXXXXXXXXXXXXXXXXX53, MXXXXXXXXXXXXXXXMXMXMXXXX, 
      MXXXXXXXXXXXXXXXXXX28, MXXXXXXXXXXXXXXXXXXXX24, 
      MXXXXXXXXXXXXXXXXXXXFXWXXX0, MXXXXXXXXXXXXXXXXXXXPXXXX, 
      MXXXXXXXXXXXXXXXXXXFXWXXX3, MXXXXXXXXXXXXXXXXXXFXWXXX4, 
      MXXXXXXXXXXXXXXXXXXFXXXXXXX0, MXXXXXXXXXXXXXXXXXXXFXWXXXXX, 
      MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, MXXXXXXXXXXXXXXXXXXFXWXXX5, 
      MXXXXXXXXXXXXXPXLXXXXXX, MXXXXXXXXXXXXXPXLXXXXXX0, 
      MXXXXXXXXXXXXXPXLXXXXXX1, MXXXXXXXXXXXXXPXLXXXXXX2, 
      MXXXXXXXXXXXXXPXLXXXXXX3, MXXXXXXXXXXXXXPXLXXXXXX4, 
      MXXXXXXXXXXXXXPXLXXXXXX5, MXXXXXXXXXXXXXPXLXXXXXX6, 
      MXXXXXXXXXXXXXPXHXXXXXX, MXXXXXXXXXXXXXPXHXXXXXX0, 
      MXXXXXXXXXXXXXPXHXXXXXX1, MXXXXXXXXXXXXXPXHXXXXXX2, 
      MXXXXXXXXXXXXXPXHXXXXXX3, MXXXXXXXXXXXXXPXHXXXXXX4, 
      MXXXXXXXXXXXXXPXHXXXXXX5, MXXXXXXXXXXXXXPXHXXXXXX6, 
      MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7, 
      MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9, 
      MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10, MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11, 
      MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12, MXXXXXXXXXXXXXXFXXXXXXXXX, 
      MXXXXXXXXXXXXXMXMPXXXXXXXX, MXXXXXXXXXXXXXPMXXXXXXX, 
      MXXXXXXXXXXXXXXXXXXXXX54, MXXXXXXXXXXXXXXXXXXXXX55, 
      MXXXXXXXXXXXXXXXXXXXXX56, MXXXXXXXXXXXXXXXXXXXXX57, 
      MXXXXXXXXXXXXXXXXXXXXX58, MXXXXXXXXXXXXXXXXXXXXX59, 
      MXXXXXXXXXXXXXXXXXXXXX60, MXXXXXXXXXXXXXXXXXXXXX61, 
      MXXXXXXXXXXXXXXXXXXXXX62, MXXXXXXXXXXXXXXXXXXXXX63, 
      MXXXXXXXXXXXXXXXXXXXXX64, MXXXXXXXXXXXXXXXXXXXXX65, 
      MXXXXXXXXXXXXXXXXXXXXX66, MXXXXXXXXXXXXXXXXXXXXX67, 
      MXXXXXXXXXXXXXXXXXXXXX68, MXXXXXXXXXXXXXXXXXXXXX69, 
      MXXXXXXXXXXXXXXXXXXXXX70, MXXXXXXXXXXXXXXXXXXXXX71, 
      MXXXXXXXXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXXXXXXXX21, 
      MXXXXXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXXXXX23, 
      MXXXXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXX8, 
      MXXXXXXXXXXXXXXFXXXXXPXXXXXXX, MXXXXXXXXXXXXXXFXXXXXPXXXXXXX0, 
      MXXXXXXXXXXXXXXFXXXXXPXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXPXXXXXXX2, 
      MXXXXXXXXXXXXXXFXXXXXPXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX1, 
      MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX3, 
      MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX4, MXXXXXXXXXXXXXXXXXX29, 
      MXXXXXXXXXXXXXXXXXXMXXXXX, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1, 
      MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2, MXXXXXXXXXXXXXXXXXXMXXX, 
      MXXXXXXXXXXXXXXXXXXMXXX0, MXXXXXXXXXXXXXXXXXXMXXX1, MXXXXXXXXXXXXXXXXXX30
      , MXXXXXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXXX, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXXX1, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXXX3, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXXX4, MXXXXXXXXXXXXXXFXXXXXXXXXXXX5, 
      MXXXXXXXXXXXXXXFXXXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXXXMXXX, 
      MXXXXXXXXXXXXXXFXXXXXXXMXXX0, MXXXXXXXXXXXXXXXXVXX, 
      MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX : std_logic;

begin
   port0o <= ( port0o0_7_port, port0o0_6_port, port0o0_5_port, port0o0_4_port, 
      port0o0_3_port, port0o0_2_port, port0o0_1_port, port0o0_0_port );
   port1o <= ( port1o0_7_port, port1o0_6_port, port1o0_5_port, port1o0_4_port, 
      port1o0_3_port, port1o0_2_port, port1o0_1_port, port1o0_0_port );
   port2o <= ( port2o0_7_port, port2o0_6_port, port2o0_5_port, port2o0_4_port, 
      port2o0_3_port, port2o0_2_port, port2o0_1_port, port2o0_0_port );
   port3o <= ( port3o0_7_port, port3o0_6_port, port3o0_5_port, port3o0_4_port, 
      port3o0_3_port, port3o0_2_port, port3o0_1_port, port3o0_0_port );
   memdatao <= ( memdatao0_7_port, memdatao0_6_port, memdatao0_5_port, 
      memdatao0_4_port, memdatao0_3_port, memdatao0_2_port, memdatao0_1_port, 
      memdatao0_0_port );
   memaddr <= ( memaddr0_15_port, memaddr0_14_port, memaddr0_13_port, 
      memaddr0_12_port, memaddr0_11_port, memaddr0_10_port, memaddr0_9_port, 
      memaddr0_8_port, memaddr0_7_port, memaddr0_6_port, memaddr0_5_port, 
      memaddr0_4_port, memaddr0_3_port, memaddr0_2_port, memaddr0_1_port, 
      memaddr0_0_port );
   ramaddr <= ( ramaddr0_7_port, ramaddr_6, ramaddr_5, ramaddr_4, ramaddr_3, 
      ramaddr_2, ramaddr_1, ramaddr_0 );
   sfrdatao <= ( sfrdatao0_7_port, sfrdatao0_6_port, sfrdatao0_5_port, 
      sfrdatao0_4_port, sfrdatao0_3_port, sfrdatao0_2_port, sfrdatao0_1_port, 
      sfrdatao0_0_port );
   sfraddr <= ( ramaddr_6, ramaddr_5, ramaddr_4, ramaddr_3, ramaddr_2, 
      ramaddr_1, ramaddr_0 );
   TraceA <= ( TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, 
      TrigOut0, TrigOut0 );
   TraceDI <= ( TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, 
      TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, 
      TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0, TrigOut0 );
   nrsto <= nrsto0;
   nrsto_nc <= nrsto_nc0;
   clkcpu_en <= clkcpu_en0;
   clkper_en <= clkper_en0;
   sfrwe <= sfrwe0;
   TrigOut <= TrigOut0;
   TraceWr <= TrigOut0;
   
   MXXXXXX : MX2 port map( A => XXXXXX8, S => XXXXXX9, B => XXXXXXXXXX6, Y => 
                           XXXXXXXXXX7);
   MXMXXXXXXXXXXXXXXXXXXXXXX : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, S => 
                           XXXXXXXXX1, B => memdatai(1), Y => 
                           MXMXXXXXXXXXXXXXXXXX);
   MXMXXXXXXXXXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, S => 
                           XXXXXXXXXX7, B => memdatai(5), Y => 
                           MXMXXXXXXXXXXXXXXXXX0);
   XXXXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => MXXXXXXXXXXXXXXXXXXXXXXX1, B =>
                           MXXXXXXXXXXXXXXXXXXXXXXX2, Y => XXXXXXXXXXXXXXXXXX);
   XXX2 : AO1B port map( A => XXXXXXXXXX8, B => XXXXXXXXXX9, C => XXXXXXXXX2, Y
                           => XXXXXX10);
   MXXXXXXXXXXXX : AO1 port map( A => MXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX, Y => MXXXXXXX4);
   XXXXXXXX1 : NOR3C port map( A => MXMPXXXXWXXX, B => XXXXXXXXXX10, C => 
                           XXXXXX11, Y => XXXXXXXXXX11);
   MXXX : OR3C port map( A => MXXXXX6, B => MXXXXXXXXXXXXXXXXLXXXXXXX0, C => 
                           MXXXXXXX4, Y => XXXXXXXXX2);
   MXMXXXXXXXXXXXXXXXXXXXX : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1, S => 
                           XXXXXXXXXX7, B => memdatai(3), Y => 
                           MXMXXXXXXXXXXXXXXX);
   MXXXX : MX2 port map( A => XXXXXX8, S => XXXXXX9, B => XXXXXXXXXX6, Y => 
                           XXXXXXXX11);
   XXXXXXXXX : OR2A port map( A => MXXXXXX1, B => XXXXXXXXXX11, Y => XXXXXX12);
   XXXXX5 : INV port map( A => XXX10, Y => XXXXXX8);
   XXXXX6 : INV port map( A => XXXXXX13, Y => XXXXXX11);
   XXXXX7 : MX2 port map( A => XXXXXX10, S => XXXXXX14, B => XXXXXX15, Y => 
                           XXXXXXX24);
   XXXXXXX3 : OR2A port map( A => MXXX16, B => XXXXXXX24, Y => XXXXXX16);
   XXXXXXX4 : MX2 port map( A => MXXXXX7, S => XXXXXX16, B => XXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0);
   XXX3 : OR3C port map( A => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX, B => 
                           MXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, Y => XXXXXX13
                           );
   XXXXX8 : OR3B port map( A => XXX11, B => XXXX17, C => XXXXXX12, Y => XXX10);
   XXXXXX2 : INV port map( A => XXXX18, Y => XXXXXXXX12);
   XXXXXX3 : INV port map( A => XXXX17, Y => XXXXXXXX13);
   XXXXXXX5 : OR3B port map( A => MXMPXXXXWXXX, B => XXXX18, C => XXXXXXXXXX12,
                           Y => XXXX17);
   XXXXXXX6 : OR3B port map( A => XXXXXXXXXXXXXX, B => XXXXXXXXXXXX3, C => 
                           XXXXXXXX14, Y => XXXXXX14);
   XXXXXX4 : XOR2 port map( A => XXXXXXXXX4, B => MXXXXXXXXXXXXXXXXXXX, Y => 
                           XXXXXXXX14);
   XXXXXXX7 : AO1C port map( A => MXXXXXXXXXXXXXXXXXXXXX1, B => MXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXXXXX, Y => XXXXXXXXX4);
   XXXXXXX8 : AO1B port map( A => MXXXXXXXXXXXXXXXXLXXXXXXX0, B => MXXXXXXX4, C
                           => XXXXXXXX14, Y => XXXXXX15);
   XXXXXXX9 : MX2A port map( A => XXX10, S => XXXXXX9, B => XXXXXXXXXX6, Y => 
                           XXXXXXXXX1);
   XXXXXXX10 : OR2B port map( A => XXXXXX13, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, Y => XXXX18);
   XXXXX9 : MX2 port map( A => XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2, S =>
                           XXXXXXXXX1, B => memdatai(2), Y => MXMXXXXXXXXXXXXX)
                           ;
   XXXXX10 : OR3B port map( A => MXXXXXX1, B => XXX11, C => XXXXXXXXXX11, Y => 
                           MXXXXXX2);
   XXXXX11 : MX2 port map( A => XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3, S 
                           => XXXXXXXXX1, B => memdatai(0), Y => 
                           MXMXXXXXXXXXXXXX0);
   XXXXX12 : OR2A port map( A => XXXX18, B => XXXXXXXXXX13, Y => XXX11);
   XXXXXXXXXX : OR3A port map( A => MXXXXX9, B => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXLXXX, C => XXXXX31, Y => 
                           XXXXX32);
   XXXXXXXXXX0 : OR3 port map( A => XFXXXXXXXXXX, B => XFXXXXXXXXXXXX, C => 
                           XXXXX33, Y => XXXXX31);
   XXXXXXX11 : OR2 port map( A => ramaddr_3, B => ramaddr_4, Y => XXXXX33);
   XXXXXXX12 : OR3 port map( A => XFXXXXXXXXXX, B => XFXXXXXXXXXXXX, C => 
                           XXXXX34, Y => XXXXX35);
   XXXXXXXXX0 : OR2 port map( A => ramaddr_3, B => ramaddr_4, Y => XXXXX34);
   XXXXX13 : OR3A port map( A => MXXXXX10, B => XXXXX35, C => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXLXXX, Y => XXXXXXX25);
   XXXXX14 : OR3A port map( A => MXXXXX10, B => XXXXX32, C => MXXXXX11, Y => 
                           XXXX19);
   XXXXXXXXXX1 : OR2 port map( A => XXXXXX17, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, Y => 
                           XXXXXXX26);
   XXX4 : MX2B port map( A => XXXXXXX26, S => MXXX17, B => XXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX);
   XXXXX15 : MX2B port map( A => MXXXX12, S => XXXX19, B => XXXXXXX27, Y => 
                           XXXXXX17);
   XXX5 : MX2B port map( A => MXXXX13, S => XXXXXXX25, B => MXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX);
   XXXXXXXXXXXXX : BUFF port map( A => nreset, Y => XXXXXXXX15);
   XXXXXXXXXXXXX0 : BUFF port map( A => nreset, Y => XXXXXXXX16);
   XXXXXXXXXXXXX1 : BUFF port map( A => nreset, Y => XXXXXXXX17);
   XXXXX16 : MX2C port map( A => MXXXX14, S => XXXXX36, B => XXXXXXXX14, Y => 
                           XFXXXXXXXXXXX);
   XXXXXXX13 : MX2C port map( A => MXXXX14, S => XXXXX36, B => XXXXXXXX14, Y =>
                           XFXXXXXXXXXXX0);
   MXMXXXXXXXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, S => 
                           XXXXXXXX11, B => memdatai(5), Y => 
                           MXMXXXXXXXXXXXXXXX0);
   MXMXXXXXXXXXXXXXXXXXXXX1 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, S => 
                           XXXXXXXX11, B => memdatai(5), Y => 
                           MXMXXXXXXXXXXXXXXX1);
   MXMXXXXXXXXXXXXXXXXXXXX2 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, S => 
                           XXXXXXXX11, B => memdatai(5), Y => 
                           MXMXXXXXXXXXXXXXXX2);
   MXMXXXXXXXXXXXXXXXXXXXX3 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3, S => 
                           XXXXXXXX11, B => memdatai(0), Y => 
                           MXMXXXXXXXXXXXXXXX3);
   MXMXXXXXXXXXXXXXXXXXXXX4 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3, S => 
                           XXXXXXXX11, B => memdatai(0), Y => 
                           MXMXXXXXXXXXXXXXXX4);
   MXMXXXXXXXXXXXXXXXXXXXX5 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1, S => 
                           XXXXXXXX11, B => memdatai(3), Y => 
                           MXMXXXXXXXXXXXXXXX5);
   MXMXXXXXXXXXXXXXXXXXXXX6 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1, S => 
                           XXXXXXXXXX7, B => memdatai(3), Y => 
                           MXMXXXXXXXXXXXXXXX6);
   MXMXXXXXXXXXXXXXXXXXXXX7 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4, S => 
                           XXXXXXXXXX7, B => memdatai(4), Y => 
                           MXMXXXXXXXXXXXXXXX7);
   MXMXXXXXXXXXXXXXXXXXXXX8 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4, S => 
                           XXXXXXXXXX7, B => memdatai(4), Y => 
                           MXMXXXXXXXXXXXXXXX8);
   MXMXXXXXXXXXXXXXXXXXXXX9 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4, S => 
                           XXXXXXXXXX7, B => memdatai(4), Y => 
                           MXMXXXXXXXXXXXXXXX9);
   MXMXXXXXXXXXXXXXXXXXXXX10 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2, S => 
                           XXXXXXXXXX7, B => memdatai(2), Y => 
                           MXMXXXXXXXXXXXXXXX10);
   MXMXXXXXXXXXXXXXXXXXXXX11 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2, S => 
                           XXXXXXXXX1, B => memdatai(2), Y => 
                           MXMXXXXXXXXXXXXXXX11);
   MXMXXXXXXXXXXXXXXXXXXXX12 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, S => 
                           XXXXXXXXX1, B => memdatai(1), Y => 
                           MXMXXXXXXXXXXXXXXX12);
   MXMXXXXXXXXXXXXXXXXXXXX13 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, S => 
                           XXXXXXXXX1, B => memdatai(1), Y => 
                           MXMXXXXXXXXXXXXXXX13);
   MXMXXXXXXXXXXXXXXXXXXXX14 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, S => 
                           XXXXXXXXX1, B => memdatai(1), Y => 
                           MXMXXXXXXXXXXXXXXX14);
   XXXXXXX14 : MX2B port map( A => MXXXXX13, S => MXXXXX14, B => XXXXXXXX18, Y 
                           => MXMXXXXXXXXXXXXXXX15);
   XXXXXXX15 : MX2B port map( A => MXXXXX13, S => MXXXXX14, B => XXXXXXXX18, Y 
                           => MXMXXXXXXXXXXXXXXX16);
   XXXXXXX16 : MX2B port map( A => MXXXXX13, S => MXXXXX14, B => XXXXXXXX18, Y 
                           => MXMXXXXXXXXXXXXXXX17);
   MXXXX0 : MX2C port map( A => XXXXXXX28, S => XXXXXXXXXX14, B => XXXXXXX29, Y
                           => MXMXXXXXXXXXXXXXXX18);
   MXXXX1 : MX2C port map( A => XXXXXXX28, S => XXXXXXXXXX14, B => XXXXXXX29, Y
                           => MXMXXXXXXXXXXXXXXX19);
   MXXXX2 : MX2C port map( A => XXXXXXX28, S => XXXXXXXXXX14, B => XXXXXXX29, Y
                           => MXMXXXXXXXXXXXXXXX20);
   XXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => MXXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, Y => XXXXXXXXXXXXXXXX0);
   XXXXXXXXXXXXXXX : OAI1 port map( A => XXXXXXXX12, B => XXXXXXXXXX13, C => 
                           MXXXXXX1, Y => XXXXXXXXXX15);
   XXXXXXXXXXXX : AO1C port map( A => MXXXXXXXXXXXXXXXXXFXXXHX, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX, C => MXMPXXXXWXXX, Y => 
                           XXXXXXXXXX13);
   XXXXXXXXXXXX0 : OR2A port map( A => XXXXXXMXXX, B => XXXXXXX25, Y => 
                           XXXXXXXXXX12);
   XXXXXXXXXXXXXXX0 : NOR2A port map( A => XXXXXXX25, B => MXXXXX12, Y => 
                           XXXXXXXXXX10);
   XXXXXXXXXXXXXXX1 : NOR3A port map( A => XXXXXXX25, B => MXXXXX12, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, Y => XXXXXXXXXX16)
                           ;
   MXXXXXXXXXX : NOR2B port map( A => MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, B => 
                           MXXX16, Y => MXXXXX15);
   MXXXXXXXXXXXX0 : OR2B port map( A => MXXXXXXXXXXXXXMXMPXXXXXX, B => MXXXXXX3
                           , Y => MXXXXXXX6);
   MXXXXXXX : OR2B port map( A => mempsacki, B => XXXXXPXXX, Y => MXXXXX16);
   MXXXXXXXXXX0 : NOR3A port map( A => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX,
                           B => MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX1, Y => MXXXXX6);
   MXXXXXXXXXX1 : NOR3C port map( A => MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, C => MXXXXX17,
                           Y => MXXXXX18);
   MXXXXXXXXXX2 : NOR2A port map( A => MXXXXX19, B => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXLXXX, Y => MXXXXX17);
   MXXXXXXXXXX3 : NOR3A port map( A => MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXX, B => 
                           XFXXXXXXXXXX0, C => XFXXXXXXXXXX1, Y => MXXXXX19);
   XXXXXXXXXXXXXXX2 : NOR3B port map( A => MXXXXXXXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXXXX17, C => XXXXXXX30, Y => XXXXXXXXXX9);
   MXXXXXXX0 : NOR3C port map( A => MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXX, Y => MXXXXX10);
   MXXXXXXX1 : NOR2B port map( A => XXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX36, Y => 
                           MXXXXX8);
   MXXXXX : NOR2 port map( A => MXXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, Y => MXXX18);
   XXXXXXXXXXXXXXXXXXX : NOR2A port map( A => XXXXXXXXXXXX4, B => 
                           XXXXXXXXXXXXXXXX0, Y => XXXXXXXXXXXXXX0);
   XXXXXXXXXXXXXXXXX : NOR2A port map( A => MXXXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX2, Y => XXXXXXXXXXXX4);
   MXXXXXXXXXXX : NOR2B port map( A => XXXXXXXX19, B => MXXXXXXXX, Y => 
                           MXXXXXX4);
   MXXXXXXXXXXXXX : NOR2A port map( A => MXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, Y => MXXXXXXXX);
   MX : NOR3A port map( A => MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX, B => 
                           XXXXXXX30, C => MXXXXXXXXXXXXXXXXLXXXXXXX1, Y => 
                           XXXXX36);
   MXXX0 : OR3C port map( A => MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, B => 
                           MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, Y => MXXXXX12)
                           ;
   MXXXXXXXXXX4 : OR3B port map( A => XXXXXXXX14, B => XXXXXXXXX2, C => 
                           XXXXXXX30, Y => MXXXXXXX7);
   XXXXXXXX2 : NOR3B port map( A => MXXXXX20, B => XXXXXXXXXX18, C => XXXXXXX25
                           , Y => XXXXXXX31);
   MXXXX3 : OR3 port map( A => MXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX2, C => MXXXXXXX8, Y => 
                           MXXXXXX6);
   MXXXXX0 : OR3A port map( A => MXXXXXXXXXXXXXXXXLXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXX0, Y => MXXXXXXX9);
   MXXX1 : AO1B port map( A => MXXX19, B => MXXXXXXX5, C => MXXXXX15, Y => 
                           MXXXXX21);
   MXXXXX1 : NOR3C port map( A => MXXXXX22, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, C => MXXX19, Y => 
                           XXXXXX18);
   XXXXXXXX3 : NOR3B port map( A => MXXXXX16, B => MXXXXX23, C => MXX5, Y => 
                           XXXXXXXXXX6);
   XXXXXXXX4 : NOR3 port map( A => XXXXXXXXXX11, B => XXXXXXXXX5, C => XXXXXX9,
                           Y => XXXXXXXXXX14);
   MXXXXX2 : NOR3B port map( A => MXXXXXXX10, B => MXXXX15, C => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, Y => 
                           MXXXXXXX11);
   XXXXXXXXXX2 : OR2A port map( A => XXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX0, Y => XXXXXXXXXX8);
   MXXXXX3 : NOR3 port map( A => MXXXXX24, B => XXXXXXX30, C => XXXXXXXXX4, Y 
                           => MXXXXXXX12);
   MXXXXX4 : NOR3A port map( A => MXXXXXXXXXXXXXXXXXXXXXXX3, B => XXXXXXX30, C 
                           => MXXXXX24, Y => XXXXXXXX20);
   XXXXXXXXXXXX1 : OR3B port map( A => MXXXXXXXXXXXXXXXXLXXXXXXX, B => 
                           XXXXXXXXXX8, C => XXXXXXX30, Y => XXXXXXXXXXXXXX);
   MXXX2 : XA1 port map( A => MXXXXX12, B => XXXXXXX32, C => MXXXXX18, Y => 
                           MXXXXX25);
   XXXXXXXXXXXX2 : NOR3A port map( A => MXXXXXXXXXXXXXXXXXXFXXXHX, B => 
                           XXXXXXXXXXXX5, C => MXXXXXXXXXXXXXXXXXFXXXHX, Y => 
                           XXXXXXXXXX18);
   XXXXXXX17 : OR3C port map( A => XXXXXXX33, B => XXXXXXX26, C => MXXX16, Y =>
                           XXXXXXXXX3);
   MXXXXXXX2 : NOR2A port map( A => MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXXX, Y => MXXXXXXX5);
   MXXXXXXX3 : NOR2A port map( A => MXXXXXXXXXXXXXXXXLXXXXXXX1, B => XXXXXXX30,
                           Y => MXXXXXXX10);
   MXXXXXXXXXX5 : NOR2A port map( A => XFXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX1, Y => MXXXXX9);
   XXXXXXXXXXXXXXXXX0 : OR2 port map( A => MXXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXX1, Y => XXXXXXXXXXXX6);
   MXXXXXXXXXXX0 : NOR2A port map( A => MXXXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX2, Y => MXXXXXX5);
   MXXXXXXXXXXXX1 : OR3A port map( A => MXXXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, Y => MXXXXXXX8);
   XXXXX17 : MX2 port map( A => MXXXXX12, S => MXXXXX25, B => XXXXXXXX21, Y => 
                           XXXXXXX27);
   MXXXX4 : AX1D port map( A => XFXXXXXXXXXX2, B => ramaddr_6, C => XXXXXXX32, 
                           Y => XXXXXXXX21);
   XXXXXXXX5 : OR3A port map( A => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX12
                           , B => MXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, Y => XXXXXXXXXX17);
   XXXXXXXXXXXXXXX3 : OR2B port map( A => XFXXXXXXXXXXXXXXXXX, B => 
                           XFXXXXXXXXXXXXXXXXX0, Y => XXXXXXXXXXXX3);
   XXXXX18 : MX2 port map( A => MXXXXXXX12, S => XXXXXXXX20, B => MXXXXX26, Y 
                           => XXXXXXX34);
   MXXXXX5 : OR2A port map( A => MXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXX1, Y => XXXXXXXX19);
   MXXX3 : AX1A port map( A => MXXXXXXXXXXXXXXXXXXX0, B => MXXX18, C => 
                           XXXXXXXXX4, Y => MXXXXX26);
   XXXXXXX18 : OR2B port map( A => MXXXXXXX4, B => XXXXXXXXXX8, Y => XXXXXXXXX6
                           );
   MXX : MX2B port map( A => XXXXXXXXX6, S => XFXXXXXXXXXXXXXXXXX0, B => 
                           XFXXXXXXXXXXXXXXXXX, Y => MXXXX14);
   XXXXX19 : MX2B port map( A => MXXXXX27, S => MXXXXX28, B => MXXXXXX7, Y => 
                           XXXXXXX33);
   MXXXXXXXXXX6 : OR2 port map( A => MXXXXXXX8, B => MXXXXXXXXXXXXXXXXXXX0, Y 
                           => MXXXXXXX13);
   MXXX4 : NOR3 port map( A => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, B => 
                           XXXXXXX25, C => MXXXXXXX11, Y => MXXXXX28);
   MXXXX5 : XO1A port map( A => XXXXXXXXX4, B => MXXXXXXX13, C => MXXXXXXXX0, Y
                           => MXXXXXX8);
   MXXXXXX0 : NOR2A port map( A => MXXXXXXXXXXXXXXXXLXXXXXXX1, B => 
                           XFXXXXXXXXXXXXXXXXX0, Y => MXXXXXXXX0);
   MXXX5 : OR2 port map( A => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, B => 
                           XXXXXXX25, Y => MXXXXX27);
   MXXXX6 : MX2 port map( A => MXXXXXX8, S => XXXXXXX34, B => MXXXX15, Y => 
                           MXXXXXX7);
   XXXXX20 : MX2 port map( A => MXXXXXX9, S => MXXXXX29, B => MXXXXXXX14, Y => 
                           XXXXXXXXX7);
   MXXX6 : OR3 port map( A => MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, B => 
                           XXXXXXX25, C => MXXXXXXX10, Y => MXXXXX29);
   MXXXX7 : AO1 port map( A => MXXXXXXX4, B => MXXXXXX6, C => 
                           XFXXXXXXXXXXXXXXXXX0, Y => MXXXXXX10);
   MXXXXXXXXXX7 : OR2 port map( A => XXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, Y => 
                           MXXXXXXX14);
   MXXXX8 : NOR2B port map( A => MXXXXXX10, B => XXXXXXXX14, Y => MXXXXXX9);
   XXXXXXXXXX3 : MX2B port map( A => MXXXXX13, S => MXXXXX14, B => XXXXXXXX18, 
                           Y => MXMXXXXXXXXXXXXX1);
   MXXX7 : MX2 port map( A => XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5, S => 
                           XXXXXXXXXX6, B => memdatai(6), Y => MXXXXX13);
   MXXX8 : XA1B port map( A => memdatai(6), B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5, C => 
                           XXXXXX9, Y => MXXXXX14);
   MXX0 : AX1D port map( A => XXXXXXXX13, B => MXXXXXX2, C => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5, Y => 
                           XXXXXXXX18);
   MXXXX9 : MX2C port map( A => MXXXXXX3, S => MXXXXX21, B => MXXXXX30, Y => 
                           MXXXXXX1);
   XXXXXXXX6 : OR2B port map( A => XXXXXXXXXX6, B => XXXXXX9, Y => XXXXXXXXXX19
                           );
   XXXXXXXX7 : XNOR2 port map( A => XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6,
                           B => memdatai(7), Y => XXXXXXXXX5);
   XXXXX21 : AX1D port map( A => XXXXXXXX13, B => XXXXXXXXXX15, C => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6, Y => 
                           XXXXXXX29);
   XXXXX22 : MX2C port map( A => memdatai(7), S => XXXXXXXXXX19, B => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6, Y => 
                           XXXXXXX28);
   MXX1 : MX2C port map( A => XXXXXXX28, S => XXXXXXXXXX14, B => XXXXXXX29, Y 
                           => MXMXXXXXXXXXXXXX2);
   XXXXXXX19 : AO1 port map( A => MXMPXXXXWXXX, B => XXXXXXXXXX16, C => 
                           MXXXXX23, Y => XXXXXX9);
   MXXX9 : AO1C port map( A => MXXXXXXX6, B => MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF
                           , C => MXX5, Y => MXXXXX23);
   MXXX10 : MX2 port map( A => MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, S => XXXXXX18,
                           B => MXXXXXXXXXXXXXMXMPXXXXXX, Y => MXXXXX30);
   MXXX11 : NOR2 port map( A => MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX, Y => MXXXXX20);
   XXXXX23 : MX2C port map( A => MXXXXXX3, S => MXXXXX21, B => MXXXXX30, Y => 
                           XXXXXXX35);
   MXXX12 : OR2 port map( A => MXXXXXXXXXXXXXMXMPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX, Y => MXXXXX22);
   MXXXX10 : MX2B port map( A => XXXXXXX24, S => XXXXXXX33, B => XXXXXXX26, Y 
                           => MXXXXXX3);
   MXX2 : AO1C port map( A => MXXXXXXXXXXXXXXXXXXX0, B => MXXXXXX4, C => 
                           MXXXXXXX4, Y => MXXXX15);
   MXXX13 : AO1A port map( A => MXXXXXX5, B => MXXXXXXXXXXXXXXXXLXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX1, Y => MXXXXX24);
   MXX3 : NOR2B port map( A => MXXXXXX6, B => MXXXXXXX4, Y => MXXXX12);
   MXXX14 : AO1 port map( A => MXXXXXXX9, B => MXXXXXXXXXXXXXXXXLXXXXXXX, C => 
                           XFXXXXXXXXXXXXXXXXX0, Y => MXXXXX11);
   MXXXX11 : OA1 port map( A => MXXXXXXXXXXXXXXXXLXXXXXXX1, B => 
                           XFXXXXXXXXXXXXXXXXX0, C => XFXXXXXXXXXXXXXXXXX, Y =>
                           XXXXXXX32);
   XXXXXXMX : MX2 port map( A => XXXXXXXX14, S => XXXXXXXXX2, B => MXXXX14, Y 
                           => XXXXXXMXXX);
   MX0 : NOR2 port map( A => MXXXXXXXXXXXXXMXMPXXXXXX, B => mempsacki, Y => 
                           MXXX16);
   MXXX15 : NOR2A port map( A => XXXXXXX33, B => XXXXXXX26, Y => MXXXXX7);
   XXXXXXXXXX4 : AO1 port map( A => XXXXXXXXXX18, B => MXXXXX12, C => 
                           XXXXXXXXXX20, Y => XXX12);
   XXXXXXXXXX5 : OR2B port map( A => mempsacki, B => XXXXXPXXX, Y => 
                           XXXXXXXXXXXX5);
   XXXXXXXX8 : NOR2 port map( A => MXXXXX20, B => XXXXXXXXXXXX5, Y => 
                           XXXXXXXXXX20);
   M : MX2B port map( A => XXX12, S => XXXXXXX31, B => MXXXX13, Y => MXX5);
   MX1 : MX2A port map( A => XXXXXXX24, S => XXXXXXXXX7, B => XXXXXXX26, Y => 
                           MXXX19);
   MX2_label : AO1 port map( A => MXXXXXXX7, B => XXXXXXXX14, C => XXXXXXX25, Y
                           => MXXX20);
   MX3 : NOR2 port map( A => MXXX20, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, Y => 
                           MXXX17);
   X : MX2B port map( A => MXXXX13, S => XXXXXXX25, B => MXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXFXXXHX0);
   MXX4 : MX2 port map( A => XXXXXXXX14, S => XXXXXXXXX2, B => MXXXX14, Y => 
                           MXXXX13);
   XXX6 : MX2C port map( A => MXXXX14, S => XXXXX36, B => XXXXXXXX14, Y => 
                           sfrdatao0_1_port);
   MXMXXXXXXXXXXXXXXXXXX : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, S => 
                           XXXXXXXXX1, B => memdatai(5), Y => MXMXXXXXXXXXXXXX3
                           );
   MXMXXXXXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4, S => 
                           XXXXXXXXX1, B => memdatai(4), Y => MXMXXXXXXXXXXXXX4
                           );
   MXMXXXXXXXXXXXXXXXXXX1 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1, S => 
                           XXXXXXXXX1, B => memdatai(3), Y => MXMXXXXXXXXXXXXX5
                           );
   MXMXXXXXXXXXXXXXXXXXX2 : MX2 port map( A => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, S => 
                           XXXXXXXXX1, B => memdatai(1), Y => MXMXXXXXXXXXXXXX6
                           );
   XXXXXXXXXXXXXXXX : OR2A port map( A => XXXXXXXX17, B => JXXXXX, Y => 
                           XXXXXXXXXXX);
   MXMWXXXXXX : NOR2A port map( A => MXMWXXXXXX0, B => XXXXXPXWX, Y => memwr);
   XXXMXMPXWXXXXXX : NOR2B port map( A => MXMWXXXXXX0, B => XXXXXPXWX, Y => 
                           dbgmempswr);
   XXXXX24 : GND port map( Y => TrigOut0);
   XXXXXXX20 : GND port map( Y => TrigOut0);
   UDRCK_inst : CLKINT port map( A => UDRCK_1, Y => UDRCK);
   UJTAG_inst : UJTAG port map( UIREG0 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX6, UIREG1
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX5, 
                           UIREG2 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX4, UIREG3
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX1, 
                           UIREG4 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX3, UIREG5
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX2, 
                           UIREG6 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, UIREG7 
                           => XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, 
                           URSTB => URSTB, UDRSH => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH, UDRCAP => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXP, UDRCK => 
                           UDRCK_1, UDRUPD => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXPX, UTDI => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, UTDO => 
                           XXXXXXXXXXXXXXXXXJXXXXX, TDI => TDI, TMS => TMS, TCK
                           => TCK, TRSTB => TRSTB, TDO => TDO);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXXXXXXX : NOR3C port map( A => 
                           MXMXXXXXXXXXXXXXXX11, B => MXMXXXXXXXXXXXXXXX2, C =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX1, B => 
                           MXMXXXXXXXXXXXXXXX9, C => MXMXXXXXXXXXXXXXXX17, Y =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXXXX : NOR3B port map( A => 
                           MXMXXXXXXXXXXXXXXX20, B => MXMXXXXXXXXXXXXXXX4, C =>
                           MXXXXXXXXXXXXXXXXXXX126, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXX27, C => MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, Y =>
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXFXXXHXX : NOR3A port map( A => XXXXXXX35, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX7, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : AO1C port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXPFF, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXX0, B => 
                           MXMXXXXXXXXXXXXXXX13, C => MXMXXXXXXXXXXXXXXX6, Y =>
                           MXXXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, B => MXXXXXXXXXXXXXXXXXX20
                           , Y => MXXXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXMXMPXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX, B => XXXXXXXXP, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX, B => 
                           MXXXXXXXXXXXXXXYXLXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX0, B => 
                           MXXXXXXXXXXXXXXYXLXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX2, B => 
                           MXXXXXXXXXXXXXXYXLXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           XXXXXXXX27, C => MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, Y =>
                           MXXXXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => XXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : XO1 port map( A => 
                           MXXXXXXXXXXXXXXYXLXXXX1, B => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXFXXXHXXXXXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, B => 
                           MXXXXXXXXXXXXXMXMPXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXX126);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXX10, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, CLK => clkcpu, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX29, Q => XXXXXXXX27);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1, CLK => clkcpu, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX29, Q => 
                           MXXXXXXXXXXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXPFFXXXXX : DFN1E0C0 port map( D => XXXXXXXXP, E 
                           => MXXXXXXXXXXXXXXXXXXXXXXX9, CLK => clkcpu, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX29, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXPFF);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXXFXWXXXXXXXXXX : OR2B port map( A 
                           => XFXXXXXXXXXX2, B => MXXXXXXXXXXXXXXXPXXXXXXXXXX, 
                           Y => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXFXWXXXXXXXXXX : OR2A port map( A =>
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX, B => XFXXXXXXXXXX2, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, B => port1o0_0_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX0 : NOR2B port map( A => 
                           port2o0_0_port, B => MXXXXXXXXXXXXXXXPXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX0);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX1 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, B => port3o0_0_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX1);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX2 : NOR3A port map( A => port1i(0), B 
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX2);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX3 : NOR3A port map( A => port3i(0), B 
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX3);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX4 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, B => port1o0_1_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX4);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX5 : NOR2B port map( A => 
                           port2o0_1_port, B => MXXXXXXXXXXXXXXXPXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX5);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX6 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, B => port3o0_1_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX6);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX7 : NOR3A port map( A => port1i(1), B 
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX7);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX8 : NOR2B port map( A => port2i(1), B 
                           => MXXXXXXXXXXXXXXXPXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX8);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX9 : NOR3A port map( A => port3i(1), B 
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX9);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX10 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, B => port1o0_2_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX10);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX11 : NOR2B port map( A => 
                           port2o0_2_port, B => MXXXXXXXXXXXXXXXPXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX11);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX12 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, B => port3o0_2_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX12);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX13 : NOR3A port map( A => port1i(2), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX13);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX14 : NOR3A port map( A => port3i(2), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX14);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX15 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, B => port1o0_3_port, C =>
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX15);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX16 : NOR2B port map( A => 
                           port2o0_3_port, B => MXXXXXXXXXXXXXXXPXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX16);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX17 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, B => port3o0_3_port, C =>
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX17);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX18 : NOR3A port map( A => port1i(3), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX18);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX19 : NOR3A port map( A => port3i(3), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX19);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX20 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, B => port1o0_4_port, C =>
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX20);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX21 : NOR2B port map( A => 
                           port2o0_4_port, B => MXXXXXXXXXXXXXXXPXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX21);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX22 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, B => port3o0_4_port, C =>
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX22);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX23 : NOR3A port map( A => port1i(4), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX23);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX24 : NOR3A port map( A => port3i(4), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX24);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX25 : NOR3A port map( A => port1i(5), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX25);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX26 : NOR2B port map( A => port2i(5), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX26);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX27 : NOR3A port map( A => port3i(5), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX27);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX28 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, B => port1o0_6_port, C =>
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX28);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX29 : NOR2B port map( A => 
                           port2o0_6_port, B => MXXXXXXXXXXXXXXXPXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX29);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX30 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXXXX0, B => port3o0_6_port, C =>
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX30);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX31 : NOR3A port map( A => port1i(6), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXMWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX31);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX32 : NOR2B port map( A => port2i(6), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX32);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX33 : NOR3A port map( A => port3i(6), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXMWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX33);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX34 : NOR3A port map( A => port1i(7), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXMWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX34);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX35 : NOR3A port map( A => port3i(7), B
                           => MXXXXXXXXXXXXXXXPXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXMWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX35);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXFXWXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXFXWXXX, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX);
   MXXXXXXXXXXXXXXXPXXXXXXXXXXMWXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXMWXXXXX, C => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1);
   MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXMWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1, B => port0o0_6_port, C 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX28, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX0 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2, B => port0i(6), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX31, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX0);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX1 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX29, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX30, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX4);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX2 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX32, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX33, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX1);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX3 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2, B => port0i(5), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX25, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX1);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX4 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1, B => port0o0_4_port, C 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX20, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX2);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX5 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2, B => port0i(4), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX23, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX3);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX6 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX0, B => port2i(4), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX24, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX4);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX7 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX21, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX22, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX5);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX3);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX8 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1, B => port0o0_3_port, C 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX15, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX6);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX9 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2, B => port0i(3), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX18, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX7);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX10 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX0, B => port2i(3), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX19, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX8);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX11 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX16, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX17, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX9);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXX0 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX2);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX12 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1, B => port0o0_2_port, C 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX10, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX10);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX13 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2, B => port0i(2), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX13, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX11);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX14 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX0, B => port2i(2), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX14, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX12);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX15 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX11, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX12, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX13);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX16 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1, B => port0o0_1_port, C 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX4, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX14);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX17 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2, B => port0i(1), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX7, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX15);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX18 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX5, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX6, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX3);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX19 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX8, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX9, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX0);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX20 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1, B => port0o0_0_port, C 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX16);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX21 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2, B => port0i(0), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX2, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX17);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX22 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX0, B => port2i(0), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX3, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX18);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX23 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX0, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX1, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX19);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXXFXWXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXFXWXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXFXWXXXXXXXX0 : NOR2A port map( A =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXXFXWXXXXXXXX0 : NOR2 port map( A =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXX29, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX2, B => XFXXXXXXXXXXXX, C
                           => MXXXXXXXXXXXXXXMWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX0);
   MXXXXXXXXXXXXXXXPXXXXXXXXXXMWXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX2, B => XFXXXXXXXXXXXX, C
                           => MXXXXXXXXXXXXXXMWXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXFXWXXXXXX0 : NOR2A port map( A => 
                           sfrwe0, B => MXXXXXXXXXXXXXXXPXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXXFXWXXXXXX : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX2, B => XFXXXXXXXXXXXX, C
                           => sfrwe0, Y => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXXFFXXXXXXXXXFXWXXXXXX0 : NOR2A port map( A => 
                           sfrwe0, B => MXXXXXXXXXXXXXXXPXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX24 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX0, B => port2i(7), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX35, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX20);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX25 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX2, B => port0i(7), C => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX34, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX21);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX36 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXX, B => port3o0_7_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX36);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX37 : NOR2B port map( A => 
                           port2o0_7_port, B => MXXXXXXXXXXXXXXXPXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX37);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX38 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXX, B => port1o0_7_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX38);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX26 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1, B => port0o0_7_port, C 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX38, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX22);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX27 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX37, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX36, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX23);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXX1 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX21, B => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX1);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXX2 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX17, B => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX18, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX0);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXX3 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX28 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX26, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX27, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX29 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX39, B => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX40, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX2);
   MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXVXXXXX30 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXX1, B => port0o0_5_port, C 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX41, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXXFXXXXXPXXXXXXXXX24);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX39 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXX, B => port3o0_5_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX40);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX40 : NOR2B port map( A => 
                           port2o0_5_port, B => MXXXXXXXXXXXXXXXPXXXXXXXXX, Y 
                           => MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX39);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXXXXXXX41 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXMWXXXXX, B => port1o0_5_port, C => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPXXXXXPXXXXXXMXXX41);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX : DFN1E1P0 port map( D => sfrdatao0_0_port, 
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           port3o0_0_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX0 : DFN1E1P0 port map( D => sfrdatao0_1_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           port3o0_1_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX1 : DFN1E1P0 port map( D => sfrdatao0_2_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           port3o0_2_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX2 : DFN1E1P0 port map( D => sfrdatao0_3_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           port3o0_3_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX3 : DFN1E1P0 port map( D => sfrdatao0_4_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           port3o0_4_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX4 : DFN1E1P0 port map( D => sfrdatao0_5_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           port3o0_5_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX5 : DFN1E1P0 port map( D => sfrdatao0_6_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           port3o0_6_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX6 : DFN1E1P0 port map( D => sfrdatao0_7_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           port3o0_7_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX7 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, CLK => clkper, PRE
                           => MXXXXXXXXXXXXXXXXXXXXX54, Q => port2o0_0_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX8 : DFN1E1P0 port map( D => sfrdatao0_1_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, CLK => clkper
                           , PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port2o0_1_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX9 : DFN1E1P0 port map( D => sfrdatao0_2_port,
                           E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, CLK => clkper
                           , PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port2o0_2_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX10 : DFN1E1P0 port map( D => sfrdatao0_3_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port2o0_3_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX11 : DFN1E1P0 port map( D => sfrdatao0_4_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port2o0_4_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX12 : DFN1E1P0 port map( D => sfrdatao0_5_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port2o0_5_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX13 : DFN1E1P0 port map( D => sfrdatao0_6_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port2o0_6_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX14 : DFN1E1P0 port map( D => sfrdatao0_7_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port2o0_7_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX15 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, CLK => clkper, PRE
                           => MXXXXXXXXXXXXXXXXXXXXX55, Q => port1o0_0_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX16 : DFN1E1P0 port map( D => sfrdatao0_1_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port1o0_1_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX17 : DFN1E1P0 port map( D => sfrdatao0_2_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port1o0_2_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX18 : DFN1E1P0 port map( D => sfrdatao0_3_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port1o0_3_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX19 : DFN1E1P0 port map( D => sfrdatao0_4_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX55, Q => 
                           port1o0_4_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX20 : DFN1E1P0 port map( D => sfrdatao0_5_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port1o0_5_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX21 : DFN1E1P0 port map( D => sfrdatao0_6_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port1o0_6_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX22 : DFN1E1P0 port map( D => sfrdatao0_7_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX0, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port1o0_7_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX23 : DFN1E1P0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, CLK => clkper, PRE 
                           => MXXXXXXXXXXXXXXXXXXXXX56, Q => port0o0_0_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX24 : DFN1E1P0 port map( D => sfrdatao0_1_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port0o0_1_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX25 : DFN1E1P0 port map( D => sfrdatao0_2_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port0o0_2_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX26 : DFN1E1P0 port map( D => sfrdatao0_3_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port0o0_3_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX27 : DFN1E1P0 port map( D => sfrdatao0_4_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port0o0_4_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX28 : DFN1E1P0 port map( D => sfrdatao0_5_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port0o0_5_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX29 : DFN1E1P0 port map( D => sfrdatao0_6_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port0o0_6_port);
   MXXXXXXXXXXXXXXXPXXXXXPXXXXXXXX30 : DFN1E1P0 port map( D => sfrdatao0_7_port
                           , E => MXXXXXXXXXXXXXXXPXXXXXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXXX56, Q => 
                           port0o0_7_port);
   MXXXXXXXXXXXXXXXXXXXXXLXMXMPXXXXXXXXXXXXX : INV port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXMXMPXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX1, B 
                           => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX2,
                           C => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXX127, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXX8, B => MXXXXXXXXXXXXXXXXXXXXX39, Y
                           => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX38, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXX127, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXXXXXX39, Y
                           => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX5)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX0 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXX1 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX40, B => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXXXX2 : NOR2B port map( A =>
                           MXXXXXXXXXXXXXXXXPXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX5, Y 
                           => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX1)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX1, B =>
                           MXXXXXXXXXXXXXXXXPXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX2, Y =>
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX1, C =>
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX3, Y 
                           => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX5, B 
                           => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXXXX4,
                           C => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0, Y =>
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX27, B => int1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX26, B => int0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXX : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXX, B => MXXXXXXXXXXXXXXXL
                           , C => MXXXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX : NOR2B port map( A => XXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXFF, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXFFXXXXX : DFN1 port map( D => XXXXXXXXXXX, CLK
                           => clk, Q => MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXFF);
   MXXXXXXXXXXXXXXXXXXXXXLXMXMPXXXXXXXXXXX : DFN1 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXX, CLK => clk, Q 
                           => MXXXXXXXXXXXXXMXMPXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXLXPMXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXXX, CLK => 
                           clk, CLR => MXXXXXXXXXXXXXXXXXXXXX54, Q => 
                           MXXXXXXXXXXXXXPMXXXXXXX);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXXX : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXXX0 : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXXXX : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXXX1 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXXX2 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXXX3 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXX : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXX0 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXX : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXX0 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXX1 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXX2 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXX3 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXXX4 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXX : OR2 port map( A => XFXXXXXXXXXXXX, B => 
                           XFXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXPMXXXXXXX);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXX0 : OR2 port map( A => ramaddr_3, B => 
                           ramaddr_4, Y => MXXXXXXXXXXXXXXXPMXXXXXXX0);
   MXXXXXXXXXXXXXXXPMXXXXX : NOR3 port map( A => MXXXXXXXXXXXXXXXPMXXXXXXX, B 
                           => MXXXXXXXXXXXXXXXPMXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXLXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXLX);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXX1 : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXX2 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXX3 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXXX4 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX2, Y => nrsto0);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX0 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX1 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX71);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX2 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX70);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX3 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX69);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX4 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX68);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX5 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX67);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX6 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX66);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX7 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX65);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX8 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX64);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX9 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX63);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX10 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX62);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX11 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX61);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX12 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX60);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX13 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX59);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX14 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX58);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX15 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX57);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX16 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX56);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX17 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX55);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX18 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX54);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX19 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX45);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX20 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX46);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX21 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX47);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX22 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX48);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX23 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX49);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX24 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX50);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX25 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX51);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX26 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX52);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX27 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX53);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX28 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX41);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX29 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX42);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX30 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX43);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX31 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX44);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX32 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX36);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX33 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX37);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXXX34 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX35);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX0 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX1 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX2 : BUFF port map( A => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX3 : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX4 : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX5 : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX6 : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX7 : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXXXX8 : BUFF port map( A => nrsto_nc0, Y => 
                           MXXXXXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXPMXXXXXXXLXXPXXXXXXXPXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXLX, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXLXXPXXXXXXXPXXXX);
   MXXXXXXXXXXXXXXXPMXXXXXXXXLXXXXXXXX : OR3C port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX3, Y => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXXLXXX);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXP : AO1B port map( A => MXXXXXXXXXXXXXXXXXXXLX, B
                           => XFXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXPPMX);
   MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXXXPXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXPPMX, B => MXXXXXXXXXXXXXPMXXXXXXX,
                           Y => MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXXXPXXXX);
   MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXXXPXXXXXXXXX : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXPPMX, B => 
                           MXXXXXXXXXXXXXXXPMXXXXXXXLXXPXXXXXXXPXXXX, C => 
                           MXXXXXXXXXXXXXPMXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXXXPXXXX);
   MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXXXXXXX : DFN1P0 port map( D => clkcpu_en0, CLK
                           => clk, PRE => MXXXXXXXXXXXXXXXXXXXXX45, Q => 
                           MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXX);
   MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXXXXXXX : DFN1P0 port map( D => clkper_en0, CLK
                           => clk, PRE => MXXXXXXXXXXXXXXXXXXXXX45, Q => 
                           MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXX);
   MXXXXXXXXXXXXXXXPMXXXXXXXXXXXX1 : DFN0 port map( D => 
                           MXXXXXXXXXXXXXMXMPXXXXXXXX, CLK => clk, Q => 
                           nrsto_nc0);
   MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXXXXX : DFN0P0 port map( D => 
                           MXXXXXXXXXXXXXXXPMXXXLXPXXXXXXXXPXXXX, CLK => clk, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => clkper_en0);
   MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXXXXX : DFN0P0 port map( D => 
                           MXXXXXXXXXXXXXXXPMXXXLXXPXXXXXXXPXXXX, CLK => clk, 
                           PRE => MXXXXXXXXXXXXXXXXXXXXX54, Q => clkcpu_en0);
   MXXXXXXXXXXXXXXXXLXXXXLXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX, B => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX, C => 
                           MXXXXXXXXXXXXXMXMPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXLXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, Y => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, Y => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXXXX0 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, Y => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, Y => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXLXMXMPXXXXXXX : INV port map( A => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2, Y => mempsacko);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXFFXXXXXXXXFXWXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXFXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXFFXXXXXXXXFXWXXX : OR3B port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX1);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXFFXXXXXXXXFXWXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, B => XFXXXXXXXXXX0, Y 
                           => MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXFFXXXXXXXXFXWX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX, C => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXFFXXXXXXXXFXWX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWXXX1, B => 
                           MXXXXXXXXXXXXXXXXXX18, Y => MXXXXXXXXXXXXXXXXXXFXWX)
                           ;
   MXXXXXXXXXXXXXXXXLXXXXLXXFXXXXXXLXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXHXXX, S => 
                           MXXXXXXXXXXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXLXXFXXXXXXLXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX2, S => 
                           MXXXXXXXXXXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXLXXFXXXXXXLXXXX1 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX3, S => 
                           MXXXXXXXXXXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXLXXFXXXXXXLXXXX2 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX4, S => 
                           MXXXXXXXXXXXXXXXXXXFXWX, B => MXXXXXXXXXXXXXXMXX, Y 
                           => MXXXXXXXXXXXXXXFXXXXXXLXXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXXFXXXXXXLXXXX3 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX5, S => 
                           MXXXXXXXXXXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXXXX : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXXXX0 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXX : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXMXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXX0 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXMXXXXXXX0, S => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXMXXXXXX : AX1B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXMXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXMXXXXXX0 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXMXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXFFXXXXXXXXFXWXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX, B => ramaddr_6, Y => 
                           MXXXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXFFXXXXXXXXFXWXXX2 : NOR2 port map( A => 
                           ramaddr_5, B => ramaddr_4, Y => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXX1 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX, S => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXX : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, C => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXLXXFXXXXXXLXXXX4 : MX2 port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX6, S => 
                           MXXXXXXXXXXXXXXXXXXFXWX, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX0, B => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXMXMPXXXX1, Y => 
                           MXXXXXXXXXXXXXMXMPXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXX2, CLK => 
                           clkper, CLR => MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXX1, CLK => 
                           clkper, CLR => MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXXXX0, CLK => 
                           clkper, CLR => MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXWXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11, E => 
                           MXXXXXXXXXXXXXXXXXXXLX, CLK => clkper, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10, E => 
                           MXXXXXXXXXXXXXXXXXXXLX, CLK => clkper, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX1);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXXXXLX, CLK => clkper, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXXXXLX, CLK => clkper, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX4);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXXXXLX, CLK => clkper, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXLXPXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, E => 
                           MXXXXXXXXXXXXXXXXXXXLX, CLK => clkper, CLR => 
                           MXXXXXXXXXXXXXXXXXXXX2, Q => MXXXXXXXXXXXXXXMXX);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX : DFN1E1P0 port map( D => sfrdatao0_0_port,
                           E => MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX, CLK => 
                           clkper, PRE => MXXXXXXXXXXXXXXXXXXXX2, Q => 
                           MXXXXXXXXXXXXXXXXXXXHXXX1);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX0 : DFN1E1C0 port map( D => XFXXXXXXXXXXX, E
                           => MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX, CLK => clkper,
                           CLR => MXXXXXXXXXXXXXXXXXXXXX35, Q => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11, E => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX, CLK => clkper, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX35, Q => 
                           MXXXXXXXXXXXXXXXXXXXHXXX);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXX : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10, E => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX, CLK => clkper, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX35, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXX0 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, E => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX, CLK => clkper, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX35, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXX1 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, E => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX, CLK => clkper, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX35, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXX2 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, E => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX, CLK => clkper, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXX35, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXXXXXXX3 : DFN1E1C0 port map( D => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, E => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXFXWX, CLK => clkper, 
                           CLR => MXXXXXXXXXXXXXXXXXXXXXXX17, Q => 
                           MXXXXXXXXXXXXXXXXLXXXXLXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX37);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXX0 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX37, C => 
                           MXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX36);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX36, B => 
                           XXXXXXXXXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => MXXXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXX : OR2 port map( A => MXXXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXX0 : OR2A port map( A => MXXXXXXXXXXXXXXXXXXXXXXXXX0,
                           B => MXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXX : OR3A port map( A => MXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXX8, C => MXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXX0 : OR3B port map( A => MXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX2, C => MXXXXXXXXXXXXXXXXXXXXX3,
                           Y => MXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXX : OR2B port map( A => MXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX3, B => MXXXXXXXXXXXXXXXXXXX2, Y
                           => MXXXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => MXXXXXXXXXXXXXXXXXXXXX5,
                           C => MXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXXXX8, Y
                           => MXXXXXXXXXXXXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXXXX8, Y
                           => MXXXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXXXX8, Y
                           => MXXXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXXXX8, Y
                           => MXXXXXXXXXXXXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX3 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXXXX8, Y
                           => MXXXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX37, B => 
                           XXXXXXXXXXXX6, Y => MXXXXXXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXX9, Y => MXXXXXXXXXXXXXXXXXXXXX12
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX9, B => MXXXXXXXXXXXXXXXXXXX10, 
                           Y => MXXXXXXXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX11, B => MXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => MXXXXXXXXXXXXXXXXXXXXX5
                           , Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX0 : OR2 port map( A => MXXXXXXX8, B 
                           => MXXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX : INV port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX : NAND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX38, Y => 
                           MXXXXXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX0 : AND2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX16, B => MXXXXXXXXXXXXXXXXXXX17,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXX);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX5, B => MXXXXXXXXXXXXXXXXXXX18, 
                           C => MXXXXXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXX20, C => MXXXXXXXXXXXXXXXXXXX21,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX3 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX18, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXXXXXX17, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX5 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXXXXX11, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX6 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX8, B => 
                           MXXXXXXXXXXXXXXXXXXX24, C => MXXXXXXXXXXXXXXXXXXX12,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX7 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX25, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX19, C => 
                           MXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXX1 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX20, C => 
                           MXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX39);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX8 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, C => MXXXXXXXXXXXXXXXXXXX,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX9);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX9 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXX28, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX10 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX29, B => MXXXXXXXXXXXXXXXXXXX30,
                           C => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX11 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXX31, A => MXXXXXXXXXXXXXXXXXXX32,
                           B => MXXXXXXXXXXXXXXXXXXXXX11, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX12 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX21, B => 
                           MXXXXXXX8, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX13 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXX33, C => MXXXXXXXXXXXXXXXXXXX11,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX14);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX14 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX34, B => MXXXXXXXXXXXXXXXXXXX35,
                           C => MXXXXXXXXXXXXXXXXXXX36, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXX2 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX38);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX0 : AO1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX39, B => MXXXXXXXXXXXXXXXXXXX40,
                           C => MXXXXXXXXXXXXXXXXXXX9, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXX41, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX15 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXX0 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX22);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXX4 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXX42, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX3 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXX43, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXX5 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX4 : AOI1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, C => XXXXXXXXXXXXXXXX0, 
                           Y => MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXX6 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, B => 
                           MXXXXXXXXXXXXXXXXXXX44, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX45, B => MXXXXXXXXXXXXXXXXXXX41,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXX : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX13);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX0 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX46, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXXXX47);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX1 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX48, B => MXXXXXXXXXXXXXXXXXXXXX,
                           C => MXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXX49);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX : OR3C port map( A => XXXXXXXXXXXXXXXX0, B 
                           => MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXXX50);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX0 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXX51, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, C => 
                           MXXXXXXXXXXXXXXXXXXX52, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX2 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX7, B => 
                           MXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX3 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXX47, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX3 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX25, C => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXX24);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX1 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX53, B => MXXXXXXXXXXXXXXXXXXX54,
                           C => MXXXXXXXXXXXXXXXXXXX55, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX4 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX56, B => MXXXXXXXXXXXXXXXXXXX57,
                           C => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX15, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX5 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX58, B => MXXXXXXXXXXXXXXXXXXX59,
                           C => MXXXXXXXXXXXXXXXXXXX60, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXX : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX1, B => 
                           XXXXXXXXXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXXXXX61);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX62, Y => MXXXXXXXXXXXXXXXXXXX63)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX0 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX64, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, C => 
                           MXXXXXXXXXXXXXXXXXXX62, Y => MXXXXXXXXXXXXXXXXXXX65)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX0 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXX42);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX2 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXX22, C => MXXXXXXXXXXXXXXXXXXX9, 
                           Y => MXXXXXXXXXXXXXXXXXXX18);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX4 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX3 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX45, B => MXXXXXXXXXXXXXXXXXXX44,
                           C => MXXXXXXXXXXXXXXXXXXPXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXX17);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX5 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, C => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Y => MXXXXXXXXXXXXXXXXXXX59
                           );
   MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX0, B => MXXXXXXXXXXXXXXXXX
                           , C => MXXXXXXXXXXXXXXLXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX2 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX44, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXXXX18, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXX15);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX4 : OR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX10, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXX66, Y => MXXXXXXXXXXXXXXXXXXX67)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX5 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXMXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, C => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => MXXXXXXXXXXXXXXXXXXX6
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX16 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX11, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX6 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX51, B => MXXXXXXXXXXXXXXXXXXX35,
                           C => MXXXXXXXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXX36);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX6 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX36, B => 
                           XXXXXXXXXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXXXXX68);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX7 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX22, B => MXXXXXXXXXXXXXXXXXXX35,
                           C => MXXXXXXXXXXXXXXXXXXXXX19, Y => 
                           MXXXXXXXXXXXXXXXXXXX19);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX1 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX64, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXX69);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXX0 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX64, B => MXXXXXXXXXXXXXXXXXXX62,
                           C => MXXXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX1, Y => MXXXXXXXXXXXXXXXXX
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX0, B => MXXXXXXXXXXXXXXXXX
                           , Y => MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX7 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => MXXXXXXXXXXXXXXXXXXX7, Y
                           => MXXXXXXXXXXXXXXXXXXX70);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX8 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX71, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX8 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX7, Y => MXXXXXXXXXXXXXXXXXXXXX17
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX9 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXX72);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX9 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX71, Y => MXXXXXXXXXXXXXXXXXXX31)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX10 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX10 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => MXXXXXXXXXXXXXXXXXXXXX2
                           , C => MXXXXXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXX60);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX11 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX33, B => MXXXXXXXXXXXXXXXXXXX73,
                           Y => MXXXXXXXXXXXXXXXXXXX20);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX11 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXXXX3, C => MXXXXXXXXXXXXXXXXXXX74
                           , Y => MXXXXXXXXXXXXXXXXXXX21);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX12 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX12 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX71, Y => MXXXXXXXXXXXXXXXXXXX75)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX13 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, B => XXXXXXXXXXXXXXXXXX,
                           C => MXXXXXXXXXXXXXXXXXXX10, Y => 
                           MXXXXXXXXXXXXXXXXXXX76);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX13 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => MXXXXXXXXXXXXXXXXXXX71, 
                           Y => MXXXXXXXXXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX14 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXXXX2, C => 
                           MXXXXXXXXXXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXXX77);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX14 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX0, B => MXXXXXXXXXXXXXXXXXXX78, 
                           Y => MXXXXXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX15 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX5, B => MXXXXXXXXXXXXXXXXXXX73
                           , Y => MXXXXXXXXXXXXXXXXXXX79);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX16 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX12, B => 
                           MXXXXXXXXXXXXXXXXXXX27, Y => MXXXXXXXXXXXXXXXXXXX80)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX22, B => MXXXXXXXXXXXXXXXXXXX78,
                           Y => MXXXXXXXXXXXXXXXXXXX81);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX0 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXX43);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXX35, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXX1 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX22, B => MXXXXXXXXXXXXXXXXXXX74,
                           Y => MXXXXXXXXXXXXXXXXXXX82);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX0 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX51, B => MXXXXXXXXXXXXXXXXXXX74,
                           Y => MXXXXXXXXXXXXXXXXXXX83);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX53, B => MXXXXXXXXXXXXXXXXXXX41,
                           Y => MXXXXXXXXXXXXXXXXXXX84);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX1 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => MXXXXXXXXXXXXXXXXXXX11,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => MXXXXXXXXXXXXXXXXXXX7, 
                           Y => MXXXXXXXXXXXXXXXXXXX85);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXX86);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX2 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX56, B => MXXXXXXXXXXXXXXXXXXX78,
                           Y => MXXXXXXXXXXXXXXXXXXX87);
   MXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX56, B => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXX88);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXX12, Y => 
                           MXXXXXXXXXXXXXXXXXXX89);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX4 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXX53, Y => MXXXXXXXXXXXXXXXXXXX90)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXX : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX53, B => MXXXXXXXXXXXXXXXXXXX2, 
                           Y => MXXXXXXXXXXXXXXXXXXX91);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXX2 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => MXXXXXXXXXXXXXXXXXXX27,
                           Y => MXXXXXXXXXXXXXXXXXXX92);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX2 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => MXXXXXXXXXXXXXXXXXXX73,
                           Y => MXXXXXXXXXXXXXXXXXXX48);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX5 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX71, B => MXXXXXXXXXXXXXXXXXXX8, 
                           Y => MXXXXXXXXXXXXXXXXXXX93);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => MXXXXXXXXXXXXXXXXXXX71,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXX0 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX7, B => MXXXXXXXXXXXXXXXXXXX8, Y
                           => MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX4
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX17 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX16, Y => 
                           MXXXXXXXXXXXXXXXXXXX45);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX1 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXX22, C => MXXXXXXXXXXXXXXXXXXX9
                           , Y => MXXXXXXXXXXXXXXXXXXX8);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX18 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX22, B => MXXXXXXXXXXXXXXXXXXX9
                           , Y => MXXXXXXXXXXXXXXXXXXX11);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX15 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXX3, Y => MXXXXXXXXXXXXXXXXXXX94);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX19 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX44, Y => MXXXXXXXXXXXXXXXXXXX22)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX20 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX44, B => MXXXXXXXXXXXXXXXXXXX3, 
                           Y => MXXXXXXXXXXXXXXXXXXX71);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX16 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX95, Y => MXXXXXXXXXXXXXXXXXXX14)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX17 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX3, B => MXXXXXXXXXXXXXXXXXXX2, Y
                           => MXXXXXXXXXXXXXXXXXXX96);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX18 : OR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX2, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX16, C => 
                           MXXXXXXXXXXXXXXXXXXX73, Y => MXXXXXXXXXXXXXXXXXXX97)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX2 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX95, B => MXXXXXXXXXXXXXXXXXXX3, 
                           Y => MXXXXXXXXXXXXXXXXXXX39);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX19 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX41, Y => MXXXXXXXXXXXXXXXXXXX34)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX21 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX41, B => MXXXXXXXXXXXXXXXXXXX3, 
                           Y => MXXXXXXXXXXXXXXXXXXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX22 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXX22, C => MXXXXXXXXXXXXXXXXXXX9
                           , Y => MXXXXXXXXXXXXXXXXXXX38);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX23 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX4, B => MXXXXXXXXXXXXXXXXXXX45
                           , Y => MXXXXXXXXXXXXXXXXXXX51);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXX98, Y => MXXXXXXXXXXXXXXXXXXX64)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX45, B => MXXXXXXXXXXXXXXXXXXX2, 
                           Y => MXXXXXXXXXXXXXXXXXXX40);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX6 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXX70, B => 
                           MXXXXXXXXXXXXXXXXXXXXX21, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX5);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX7 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX74, B => MXXXXXXXXXXXXXXXXXXX56,
                           C => MXXXXXXXXXXXXXXXXXXX76, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX8 : NOR3C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX6, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX38, C => 
                           MXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX9 : OA1A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX4, B => MXXXXXXXXXXXXXXXXXXXXX5,
                           C => MXXXXXXXXXXXXXXXXXXX5, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX7);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX10 : OAI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX74, B => MXXXXXXXXXXXXXXXXXXX0, 
                           C => MXXXXXXXXXXXXXXXXXXX79, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX8);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX11 : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX9);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX3 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX81, B => MXXXXXXXXXXXXXXXXXXX80,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXVXX1);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX20 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX21 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX3, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Y => MXXXXXXXXXXXXXXXXXXX98
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX22 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXX44);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX23 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, Y => 
                           MXXXXXXXXXXXXXXXXXXX41);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXX3 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Y => MXXXXXXXXXXXXXXXXXXX95
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX24 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXX99, Y => MXXXXXXXXXXXXXXXXXXX46)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX25 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX100, B => MXXXXXXXXXXXXXXXXXXX94
                           , Y => MXXXXXXXXXXXXXXXXXXX23);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX24 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, B => 
                           MXXXXXXXXXXXXXXXXXXX3, Y => MXXXXXXXXXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX25 : AO1B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX16, B => 
                           MXXXXXXXXXXXXXXXXXXX14, C => MXXXXXXXXXXXXXXXXXXX97,
                           Y => MXXXXXXXXXXXXXXXXXXX12);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX26 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXX23, C => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Y => MXXXXXXXXXXXXXXXXXXX33
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXMX : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX23, S => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Y => MXXXXXXXXXXXXXXXXXXX1)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX26 : OA1A port map( A => XXXXXXXXXXXX6, 
                           B => MXXXXXXXXXXXXXXXXXXX96, C => 
                           MXXXXXXXXXXXXXXXXXXX48, Y => MXXXXXXXXXXXXXXXXXXX16)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX27 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX74, B => MXXXXXXXXXXXXXXXXXXX66,
                           C => MXXXXXXXXXXXXXXXXXXX47, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX27 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX16, B => MXXXXXXXXXXXXXXXXXXX3
                           , Y => MXXXXXXXXXXXXXXXXXXX99);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX28 : NOR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXXX45, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXX26);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX4 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX10, B => XXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXX34, Y => MXXXXXXXXXXXXXXXXXXX101
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX5 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXXX64, C => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXX102);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX29 : OR3B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX11, C => MXXXXXXXXXXXXXXXXXXX2, 
                           Y => MXXXXXXXXXXXXXXXXXXX58);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX28 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXXX98, C => 
                           MXXXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXXX56);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX6 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX98, B => 
                           MXXXXXXXXXXXXXXXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXXX74, Y => MXXXXXXXXXXXXXXXXXXX103
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXX4 : OR2A port map( A => XXXXXXXXXXXX6
                           , B => MXXXXXXXXXXXXXXXXXXX40, Y => 
                           MXXXXXXXXXXXXXXXXXXX104);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX7 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX40, B => MXXXXXXXXXXXXXXXXXXX74,
                           Y => MXXXXXXXXXXXXXXXXXXX105);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX8 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX10, B => XXXXXXXXXXXX6, C => 
                           MXXXXXXXXXXXXXXXXXXX106, Y => 
                           MXXXXXXXXXXXXXXXXXXX107);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXX5 : XNOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX23, B => 
                           MXXXXXXXXXXXXXXXXXXXXX4, Y => 
                           MXXXXXXXXXXXXXXXXXXX108);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXX1 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX2, Y => MXXXXXXXXXXXXXXXXXXX106)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX29 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXXXXXX3, C => MXXXXXXXXXXXXXXXXXXX2,
                           Y => MXXXXXXXXXXXXXXXXXXX66);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX6 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX106, B => MXXXXXXXXXXXXXXXXXXX8,
                           Y => MXXXXXXXXXXXXXXXXXXX109);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX30 : OR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX24, B => MXXXXXXXXXXXXXXXXXXX2
                           , C => MXXXXXXXXXXXXXXXXXXX73, Y => 
                           MXXXXXXXXXXXXXXXXXXX29);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX30 : OA1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXX31, Y => MXXXXXXXXXXXXXXXXXXX110
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX31 : OA1B port map( C => 
                           MXXXXXXXXXXXXXXXXXXX49, A => MXXXXXXXXXXXXXXXXXXX71,
                           B => MXXXXXXXXXXXXXXXXXXX38, Y => 
                           MXXXXXXXXXXXXXXXXXXX111);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX12 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX14, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, C => 
                           MXXXXXXXXXXXXXXXXXXX112, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX10);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX13 : AO1D port map( A => 
                           MXXXXXXXXXXXXXXXXXXX32, B => MXXXXXXXXXXXXXXXXXXX74,
                           C => MXXXXXXXXXXXXXXXXXXX113, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX11);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX31 : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX98, B => 
                           MXXXXXXXXXXXXXXXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXXX38, Y => MXXXXXXXXXXXXXXXXXXX113
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX17 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX19, B => XXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX16);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX32 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX114, Y => MXXXXXXXXXXXXXXXXXXX57
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX9 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX22, B => XXXXXXXXXXXX6, Y => 
                           MXXXXXXXXXXXXXXXXXXX62);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX3 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX10, Y => MXXXXXXXXXXXXXXXXXXX52)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX33 : OA1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXX22, C => 
                           MXXXXXXXXXXXXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXX114);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX34 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX9, B => MXXXXXXXXXXXXXXXXXXX10, 
                           Y => MXXXXXXXXXXXXXXXXXXX73);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX14 : AOI1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX41, B => 
                           MXXXXXXXXXXXXXXXXXXXXX25, C => 
                           MXXXXXXXXXXXXXXXXXXX112, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX4);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX32 : OR2B port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXX66, Y => MXXXXXXXXXXXXXXXXXXX115
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX25);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX35 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXX98, C => 
                           MXXXXXXXXXXXXXXXXXXXXX24, Y => 
                           MXXXXXXXXXXXXXXXXXXX112);
   MXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX98, B => 
                           MXXXXXXXXXXXXXXXXXXXXX24, C => 
                           MXXXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX4 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXX8, Y => MXXXXXXXXXXXXXXXXXXX54);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX4 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX26, B => MXXXXXXXXXXXXXXXXXXX0
                           , Y => MXXXXXXXXXXXXXXXXXXX55);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX7 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXXX78, Y => MXXXXXXXXXXXXXXXXXXX116
                           );
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX5 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX45, B => MXXXXXXXXXXXXXXXXXXX78,
                           Y => MXXXXXXXXXXXXXXXXXXX53);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX33 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX19, B => MXXXXXXX8, Y => 
                           MXXXXXXXXXXXXXXXXXXX78);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX36 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX37, B => 
                           XXXXXXXXXXXX6, Y => MXXXXXXXXXXXXXXXXXXX74);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX10 : NOR2 port map( A => MXXXXXXX8
                           , B => MXXXXXXXXXXXXXXXXXXX34, Y => 
                           MXXXXXXXXXXXXXXXXXXX117);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX37 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXXXXXXXX26, Y => MXXXXXXXXXXXXXXXXXXX9
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXMX0 : MX2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX24, S => 
                           MXXXXXXXXXXXXXXXXXXXXX4, B => 
                           MXXXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXMXXX);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX38 : AO1C port map( A => 
                           MXXXXXXXXXXXXXXXXXXX96, B => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX0, C => 
                           MXXXXXXXXXXXXXXXXXXX37, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX5);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX8 : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX96, B => MXXXXXXXXXXXXXXXXXXX78,
                           Y => MXXXXXXXXXXXXXXXXXXX118);
   MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXX1 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, B => 
                           MXXXXXXXXXXXXXXXXXXX96, Y => MXXXXXXXXXXXXXXXXXXX119
                           );
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXX11 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX11, B => MXXXXXXXXXXXXXXXXXXX96,
                           Y => MXXXXXXXXXXXXXXXXXXXXXXXVXXXX6);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX39 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX26, B => 
                           MXXXXXXXXXXXXXXXXXXX96, Y => MXXXXXXXXXXXXXXXXXXX37)
                           ;
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX0 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX1 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX0, B => MXXXXXXXXXXXXXXXXXXXXXX
                           , Y => MXXXXXXXXXXXXXXLXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX2 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXX1, B => MXXXXXXXXXXXXXXXXXXXXXX
                           , Y => MXXXXXXXXXXXXXXLXXXXXXXXXXXX2);
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXXXX3 : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX28, B => 
                           MXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXXXX3);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX40 : AO1 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXXXXXXXX26, Y => MXXXXXXXXXXXXXXXXXXX4
                           );
   MXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX : OR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX51, B => MXXXXXXXXXXXXXXXXXXX39,
                           Y => MXXXXXXXXXXXXXXXXXXX120);
   MXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX : AO1 port map( A => MXXXXXXXXXXXXXXXXXXX120
                           , B => MXXXXXXXXXXXXXXXXXXXXX26, C => 
                           MXXXXXXXXXXXXXXXXXXX121, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXVXX);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXX : NOR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXX120, B => MXXXXXXXXXXXXXXXXXXX73
                           , Y => MXXXXXXXXXXXXXXXXXXX122);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXX6 : OR2B port map( A => XXXXXXXXXXXX6
                           , B => MXXXXXXXXXXXXXXXXXXX39, Y => 
                           MXXXXXXXXXXXXXXXXXXX123);
   MXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX : NOR3 port map( A => 
                           MXXXXXXXXXXXXXXXXXXX98, B => 
                           MXXXXXXXXXXXXXXXXXXXXX24, C => MXXXXXXXXXXXXXXXXXXX8
                           , Y => MXXXXXXXXXXXXXXXXXXX121);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX34 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX22, B => 
                           MXXXXXXXXXXXXXXXXXXXXX26, Y => 
                           MXXXXXXXXXXXXXXXXXXX35);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX41 : OR2A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX19, B => 
                           MXXXXXXXXXXXXXXXXXXXXX22, Y => 
                           MXXXXXXXXXXXXXXXXXXX10);
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXX42 : NOR2 port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX27, B => 
                           MXXXXXXXXXXXXXXXXXXX23, Y => MXXXXXXXXXXXXXXXXXXX32)
                           ;
   MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXX35 : NOR3A port map( A => 
                           MXXXXXXXXXXXXXXXXXXXXX24, B => 
                           MXXXXXXXXXXXXXXXXXXXXX3, C => 
                           MXXXXXXXXXXXXXXXXXXXXX23, Y => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX27);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXXXX, CLK => clkper, CLR => 
                           MXXXXXXXXXXXXXXXXXXXXX29, Q => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXX30, CLK => clkper, CLR => 
                           nrsto0, Q => MXXXXXXXXXXXXXXXXXXXXXX0);
   MXXXXXXXXXXXXXXLXXXVXXXXXXX : DFN1C0 port map( D => MXXXXXXXXXXXXXXXXXXXXXX,
                           CLK => clkper, CLR => nrsto0, Q => 
                           MXXXXXXXXXXXXXXLXXXVXX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXX0, CLK => clkper, CLR => 
                           nrsto0, Q => MXXXXXXXXXXXXXXXXXXXXXX);
   MXXXXXXXXXXXXXXLXXXVXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX, CLK => clkper, 
                           CLR => nrsto0, Q => MXXXXXXXXXXXXXXLXXXVX);
   MXXXXXXXXXXXXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXXXX, CLK => clkper, 
                           CLR => nrsto0, Q => MXXXXXXXXXXXXXXXXXXXXX30);
   MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXXXXXXX0, CLK => clkper, 
                           CLR => nrsto0, Q => MXXXXXXXXXXXXXXXXXXXXXXXXLXX);
   MXXXXXXXXXXXXXXLXXXVXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX, CLK => clkper, CLR => 
                           nrsto0, Q => MXXXXXXXXXXXXXXLXXXVX0);
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXX : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXXXX0, CLK => clkper, CLR =>
                           nrsto0, Q => MXXXXXXXXXXXXXXLXXXXXXXXXX);
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXX0 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXXXX1, CLK => clkper, CLR =>
                           nrsto0, Q => MXXXXXXXXXXXXXXLXXXXXXXXXX1);
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXX1 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXXXX2, CLK => clkper, CLR =>
                           nrsto0, Q => MXXXXXXXXXXXXXXLXXXXXXXXXX2);
   MXXXXXXXXXXXXXXLXXXXXXXXXXXXXXX2 : DFN1C0 port map( D => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXXXX3, CLK => clkper, CLR =>
                           nrsto0, Q => MXXXXXXXXXXXXXXLXXXXXXXXXX0);
   MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX : NOR2B port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX1, B => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX, Y => MXXXXXXXXXXXXXXXX1)
                           ;
   MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX0 : XOR2 port map( A => MXXXXXXXXXXXXXXXX2, 
                           B => MXXXXXXXXXXXXXXLXXXXXXXXXX0, Y => 
                           MXXXXXXXXXXXXXXXXXXXXX28);
   MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXXX1 : AND3 port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX1, C => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX2, Y => MXXXXXXXXXXXXXXXX2
                           );
   MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX0 : XOR2 port map( A => MXXXXXXXXXXXXXXXX1, B
                           => MXXXXXXXXXXXXXXLXXXXXXXXXX2, Y => 
                           MXXXXXXXXXXXXXXXXXXXX1);
   MXXXXXXXXXXXXXXXXXXLXXXXXXXXXXX1 : XOR2 port map( A => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX, B => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX1, Y => 
                           MXXXXXXXXXXXXXXXXXXXX0);
   XXXYXXXXXX : XYXX0008 port map( XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX => 
                           UDRCK, XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXX0 => 
                           URSTB, XXXXXXXXXXXXXXXXXJXXXXX => 
                           XXXXXXXXXXXXXXXXXJXXXXX, XLX => clk, XXXXXXXX => 
                           XXXXXXXX17, JXXXXX => JXXXXX, XXXXXX => AuxOut, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXX, XXXXXXXX0 
                           => XXXXXXXX26, MXMXXXXXXXX => memdatao0_5_port, 
                           MXMXXXX(15) => memaddr0_15_port, MXMXXXX(14) => 
                           memaddr0_14_port, MXMXXXX(13) => memaddr0_13_port, 
                           MXMXXXX(12) => memaddr0_12_port, MXMXXXX(11) => 
                           memaddr0_11_port, MXMXXXX(10) => memaddr0_10_port, 
                           MXMXXXX(9) => memaddr0_9_port, MXMXXXX(8) => 
                           memaddr0_8_port, MXMXXXX(7) => memaddr0_7_port, 
                           MXMXXXX(6) => memaddr0_6_port, MXMXXXX(5) => 
                           memaddr0_5_port, MXMXXXX(4) => memaddr0_4_port, 
                           MXMXXXX(3) => memaddr0_3_port, MXMXXXX(2) => 
                           memaddr0_2_port, MXMXXXX(1) => memaddr0_1_port, 
                           MXMXXXX(0) => memaddr0_0_port, XXXXXXX(19) => 
                           TraceDO(19), XXXXXXX(18) => TraceDO(18), XXXXXXX(17)
                           => TraceDO(17), XXXXXXX(16) => TraceDO(16), 
                           XXXXXXX(15) => TraceDO(15), XXXXXXX(14) => 
                           TraceDO(14), XXXXXXX(13) => TraceDO(13), XXXXXXX(12)
                           => TraceDO(12), XXXXXXX(11) => TraceDO(11), 
                           XXXXXXX(10) => TraceDO(10), XXXXXXX(9) => TraceDO(9)
                           , XXXXXXX(8) => TraceDO(8), XXXXXXX(7) => TraceDO(7)
                           , XXXXXXX(6) => TraceDO(6), XXXXXXX(5) => TraceDO(5)
                           , XXXXXXX(4) => TraceDO(4), XXXXXXX(3) => TraceDO(3)
                           , XXXXXXX(2) => TraceDO(2), XXXXXXX(1) => TraceDO(1)
                           , XXXXXXX(0) => TraceDO(0), 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX6, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXPX => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXPX, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX3, 
                           XXXXXXXX1 => XXXXXXXX27, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXP => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXP, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXH, 
                           MXMXXXX0(3) => membank(3), MXMXXXX0(2) => membank(2)
                           , MXMXXXX0(1) => membank(1), MXMXXXX0(0) => 
                           membank(0), MXMXXXXXXXX0 => memdatao0_7_port, 
                           XXXXXXXX2 => XXXXXXXX22, MXMXXXXXXXX1 => 
                           memdatao0_3_port, MXMXXXXXXXX2 => memdatao0_0_port, 
                           XXXXXXXX3 => XXXXXXXX23, XXXXXXXX4 => XXXXXXXX24, 
                           XXXXXXXX5 => XXXXXXXX25, XXXXXXXXP => XXXXXXXXP, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX1 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX2, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX2 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX4, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX3 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX5, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX4 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX5 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX0, 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX6 => 
                           XXXXXXXXXXXXXXXXXXPXXXJXXXXPXXXXXXXXXXXXXXX1, 
                           XXXXXX0 => nreset, 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6, 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0 => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5, 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1 => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX0, 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2 => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4, 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3 => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX1, 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX4 => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX2, 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX5 => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX, 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX6 => 
                           XXXXXXXXXXXXXXXXXXHXLXXXXXXXXXXXPXXXXXXXX3, 
                           XXXXXXXX6 => XXXXXXXX15, XXXXXXXX7 => XXXXXXXX16, 
                           XXXXXPXWX => XXXXXPXWX, XXXXXPXXX => XXXXXPXXX, 
                           XXXXXXXX8 => BreakOut, XXXXXXX0 => BreakIn, XXXXXXX1
                           => XXXXXXX35, MXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXX6, MXMPXXXXX => mempsacki);
   XXXYXXXXXX0 : XYXX0007 port map( XLXXPX => clkcpu, MXXXXXXXXXXXXXXXXXXXXXXXX
                           => MXXXXXXXXXXXXXXXXXXXXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXX => 
                           MXMXXXXXXXXXXXXX3, MXMXXXXXXXXXXXXXXX => 
                           MXMXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXPXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXFXXXHX => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX, 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, MXXXXXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXYXLXXXXXX
                           => MXXXXXXXXXXXXXXYXLXXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX18, 
                           MXXXXXXXXXXXXXXYXLXXXXXX0 => 
                           MXXXXXXXXXXXXXXYXLXXXXXX0, MXXXXXXXXXXXXXXYXLXXXXXX1
                           => MXXXXXXXXXXXXXXYXLXXXXXX, MXXXXXXXXXXXXXXXXPPMX 
                           => MXXXXXXXXXXXXXXXXPPMX, 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, MXXXXXXXXXXXXXXYXXXXXX 
                           => MXXXXXXXXXXXXXXYXXXXXX, MXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXXXXXXXX1 
                           => MXXXXXXXXXXXXXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXX3
                           => MXXXXXXXXXXXXXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXXXX5
                           => MXXXXXXXXXXXXXXXXXXXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX13, 
                           MXXXXXXXXXXXXXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, 
                           MXXXXXXXXXXXXXXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX19, 
                           MXXXXXXXXXXXXXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX16, 
                           MXXXXXXXXXXXXXXXXXXXXXXX10 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXXXXXXXXXX11 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXXX0 
                           => MXXXXXXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXMWXXXXXXX
                           => MXXXXXXXXXXXXXXMWXXXXXXX0, 
                           MXXXXXXXXXXXXXXMWXXXXXXX0 => 
                           MXXXXXXXXXXXXXXMWXXXXXXX, MXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXX126, MXXXXXXXXXXXXXXXXXXLLXX => 
                           MXXXXXXXXXXXXXXXXXXLLXX, MXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXYXXXX => 
                           MXXXXXXXXXXXXXXYXXXX, MXXXXXXXXXXXXXXYXXXX0 => 
                           MXXXXXXXXXXXXXXYXXXX0, MXXXXXXXXXXXXXXYXXXX1 => 
                           MXXXXXXXXXXXXXXYXXXX2, MXXXXXXXXXXXXXXXXXFXXXHX => 
                           MXXXXXXXXXXXXXXXXXFXXXHX, MXXXXXXXXXXXXXXYXLXXXX => 
                           MXXXXXXXXXXXXXXYXLXXXX0, MXXXXXXXXXXXXXXXXXXPXXXXXX 
                           => MXXXXXXXXXXXXXXXXXXPXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, MXMXXXXXXXXXXXXXXX0 
                           => MXMXXXXXXXXXXXXXXX20, MXMXXXXXXXXXXXXXXX1 => 
                           MXMXXXXXXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX, 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, MXMXXXXXXXXXXXXXXX2 =>
                           MXMXXXXXXXXXXXXXXX17, MXMXXXXXXXXXXXXXXX3 => 
                           MXMXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXMXMPXXXXXXX => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, 
                           MXMXXXXXXXXXXXXXXX4 => MXMXXXXXXXXXXXXXXX14, 
                           MXMXXXXXXXXXXXXXXX5 => MXMXXXXXXXXXXXXXXX4, 
                           MXMXXXXXXXXXXXXXXX6 => MXMXXXXXXXXXXXXXXX2, 
                           MXMXXXXXXXXXXXXXXX7 => MXMXXXXXXXXXXXXXXX11, 
                           MXMXXXXXXXXXXXXXXXXX => MXMXXXXXXXXXXXXXXXXX0, 
                           MXMXXXXXXXXXXXXXXXXX0 => MXMXXXXXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX, MXMXXXXXXXXXXXXXXX8 => 
                           MXMXXXXXXXXXXXXXXX13, MXMXXXXXXXXXXXXXXX9 => 
                           MXMXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXX10, XXXXXXXXXXXXXXXXXX => 
                           XXXXXXXXXXXXXXXXXX, MXVX => movx, 
                           MXMXXXXXXXXXXXXXXX10 => MXMXXXXXXXXXXXXXXX16, 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, 
                           MXMXXXXXXXXXXXXXXX11 => MXMXXXXXXXXXXXXXXX10, 
                           MXMXXXXXXXXXXXXXXX12 => MXMXXXXXXXXXXXXXXX19, 
                           MXMXXXXXXXXXXXXXXX13 => MXMXXXXXXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX, 
                           MXMXXXXXXXXXXXXXXX14 => MXMXXXXXXXXXXXXXXX5, 
                           MXMXXXXXXXXXXXXXXX15 => MXMXXXXXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXYXLXXXX0 => MXXXXXXXXXXXXXXYXLXXXX2, 
                           MXXXXXXXXXXXXXXYXX => MXXXXXXXXXXXXXXYXX1, 
                           MXMXXXXXXXXXXXXXXX16 => MXMXXXXXXXXXXXXXXX0, 
                           MXMXXXXXXXXXXXXXXX17 => MXMXXXXXXXXXXXXXXX18, 
                           MXXXXXXXXXXXXXXYXLXXXX1 => MXXXXXXXXXXXXXXYXLXXXX1, 
                           MXXXXXXXXXXXXXXYXLXXXX2 => MXXXXXXXXXXXXXXYXLXXXX, 
                           MXXXXXXXXXXXXXXYXX0 => MXXXXXXXXXXXXXXYXX0, 
                           MXXXXXXXXXXXXXXYXXXX2 => MXXXXXXXXXXXXXXYXXXX1, 
                           MXXXXXXXXXXXXXXYXX1 => MXXXXXXXXXXXXXXYXX, 
                           MXMXXXXXXXXXXXXXXX18 => MXMXXXXXXXXXXXXXXX15, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX, MXXXXXXXXXXXXXXXXYXLXXXXX
                           => MXXXXXXXXXXXXXXXXYXLXXXXX, MXMXXXXXXXXXXXXXXX19 
                           => MXMXXXXXXXXXXXXXXX7, MXMXXXXXXXXXXXXXXX20 => 
                           MXMXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXPXXLXX => 
                           MXXXXXXXXXXXXXXXXXXPXXLXX, 
                           MXXXXXXXXXXXXXXXXXMXVXWXXX => 
                           MXXXXXXXXXXXXXXXXXMXVXWXXX, MXXXXXXXXXXXXXXXXXXX1 =>
                           MXXXXXXXXXXXXXXXXXXX105, MXXXXXXXXXXXXXXXXXXLL => 
                           MXXXXXXXXXXXXXXXXXXLL, XXXXXXXX => XXXXXXXX27, 
                           MXXXXXXXXXXXXXXXXXXXXXPFF => 
                           MXXXXXXXXXXXXXXXXXXXXXPFF, MXMXXXXXXXXXXXXX0 => 
                           MXMXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXX21, MXMXXXXXXXXXXXXX1 => 
                           MXMXXXXXXXXXXXXX6, MXMXXXXXXXXXXXXX2 => 
                           MXMXXXXXXXXXXXXX, MXMXXXXXXXXXXXXX3 => 
                           MXMXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXX4 => 
                           MXMXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXX5 => 
                           MXMXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXX6 => 
                           MXMXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXMXMPXXXXX => 
                           MXXXXXXXXXXXXXMXMPXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, MXXXXXXXXXXXXXXXXXXX2
                           => MXXXXXXXXXXXXXXXXXXX125, MXXXXXXXXXXXXXXXXXXX3 =>
                           MXXXXXXXXXXXXXXXXXXX124, MXXXXXXXXXXXXXXMWXXXXX => 
                           MXXXXXXXXXXXXXXMWXXXXX, MXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXX37, MXXXXXXXXXXXXXXXXYXLXXXXX0
                           => MXXXXXXXXXXXXXXXXYXLXXXXX2, 
                           MXXXXXXXXXXXXXXXXYXLXXXXX1 => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX1, 
                           MXXXXXXXXXXXXXXXXYXLXXXXX2 => 
                           MXXXXXXXXXXXXXXXXYXLXXXXX0, MXXXXXXXXXXXXXXXXXXXXX0 
                           => MXXXXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXXXXXXXX1
                           => MXXXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXXX2
                           => MXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXX3 
                           => MXXXXXXXXXXXXXXXXXXXXX36, MXXXXXXXXXXXXXXXXXXXXX4
                           => MXXXXXXXXXXXXXXXXXXXXX26, MXXXXXXXXXXXXXXXXXXXXX5
                           => MXXXXXXXXXXXXXXXXXXXXX23, MXXXXXXXXXXXXXXXXXXXXX6
                           => MXXXXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXXXX7 
                           => MXXXXXXXXXXXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXXXXXX8
                           => MXXXXXXXXXXXXXXXXXXXXX3);
   XXXYXXXXXX1 : XYXX0006 port map( MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, XLXPXX => clkper, 
                           MXXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXXX18, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX2, XFXXXXXXXXXX => 
                           XFXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXPXWXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, 
                           MXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXX23, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXXXX
                           => MXXXXXXXXXXXXXXXXXXXXX40, 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, MXXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXXX105, MXXXXXXXXXXXXXXXXXXXXX0 
                           => MXXXXXXXXXXXXXXXXXXXXX39, MXXXXXXXXXXXXXXYXXXX =>
                           MXXXXXXXXXXXXXXYXXXX1, MXXXXXXXXXXXXXXYXXXX0 => 
                           MXXXXXXXXXXXXXXYXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6, 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX, 
                           MXXXXXXXXXXXXXXXXVXXXXXX => MXXXXXXXXXXXXXXXXVXXXXXX
                           , MXXXXXXXXXXXXXXXXVXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXFX => 
                           MXXXXXXXXXXXXXXFX0, MXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXX125, MXXXXXXXXXXXXXXXXVXXXXXX1 
                           => MXXXXXXXXXXXXXXXXVXXXXXX1, MXXXXXXXXXXXXXXXXXX =>
                           MXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXX27, MXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXL => 
                           MXXXXXXXXXXXXXXXL, MXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXX124, MXXXXXXXXXXXXXXFX0 => 
                           MXXXXXXXXXXXXXXFX, MXXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXX38, MXXXXXXXXXXXXXXXXVXXXXXX2 
                           => MXXXXXXXXXXXXXXXXVXXXXXX3, 
                           MXXXXXXXXXXXXXXXXVXXXXXX3 => 
                           MXXXXXXXXXXXXXXXXVXXXXXX2, MXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXX26, MXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXFXXXXX => 
                           MXXXXXXXXXXXXXXXXXXFXXXXX, MXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXX25, MXXXXXXXXXXXXXXXXPXXXXXXXX0 
                           => MXXXXXXXXXXXXXXXXPXXXXXXXX1, 
                           MXXXXXXXXXXXXXXFXWXXX => MXXXXXXXXXXXXXXFXWXXX, 
                           MXXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXXX127, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXX3 =>
                           MXXXXXXXXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXPXXXXXXXX1 
                           => MXXXXXXXXXXXXXXXXPXXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXPXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX9, XXMXXXXXXX => ramaddr_4
                           , MXXXXXXXXXXXXXXXXXX4 => MXXXXXXXXXXXXXXXXXX23, 
                           XXXXX => int0a, MXXXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXX36, XXXXX0 => int1a, XXXX => 
                           int2, XXXX0 => int3, XXXX1 => int4, XXXX2 => int5, 
                           XXXX3 => int6, XXXX4 => int7, 
                           MXXXXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXXXXX44,
                           MXXXXXXXXXXXXXXXXXXXX1 => MXXXXXXXXXXXXXXXXXXXX22, 
                           MXXXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXXXX21, 
                           MXXXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXXXX20, 
                           MXXXXXXXXXXXXXXXXXXXX4 => MXXXXXXXXXXXXXXXXXXXX19, 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX => 
                           MXXXXXXXXXXXXXXXXXFXXXHXXX, MXXXXXXXXXXXXXXXXXFXXXHX
                           => MXXXXXXXXXXXXXXXXXFXXXHX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, XFXXXXXX(7) => 
                           sfrdatao0_7_port, XFXXXXXX(6) => sfrdatao0_6_port, 
                           XFXXXXXX(5) => sfrdatao0_5_port, XFXXXXXX(4) => 
                           sfrdatao0_4_port, XFXXXXXX(3) => sfrdatao0_3_port, 
                           XFXXXXXX(2) => sfrdatao0_2_port, XFXXXXXX(1) => 
                           sfrdatao0_1_port, XFXXXXXX(0) => sfrdatao0_0_port, 
                           XFXXXXXXXXXXX => XFXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXXXXXXXX4 => MXXXXXXXXXXXXXXXXXXXXX43,
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXXXXXXXX5 => MXXXXXXXXXXXXXXXXXXXXX42,
                           MXXXXXXXXXXXXXXXXXXXXX6 => MXXXXXXXXXXXXXXXXXXXXX41)
                           ;
   XXXYXXXXXX2 : XYXX0005 port map( MXXXXXXXXXXXXXXYXLXXXXXX => 
                           MXXXXXXXXXXXXXXYXLXXXXXX1, MXXXXXXXXXXXXXXYXLXXXXXX0
                           => MXXXXXXXXXXXXXXYXLXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXXXXX2,
                           MXXXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXXXX1
                           , MXXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXXXXXXX1 => MXXXXXXXXXXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXXXX12, 
                           MXXXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXXXX13, 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX, MXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1, 
                           MXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX4, 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX, XFXXXXXXXXXX => 
                           XFXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0 => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1, XXXX => int1, 
                           MXXXXXXXXXXXXXXXX1 => MXXXXXXXXXXXXXXXX8, XXXX0 => 
                           int0, MXXXXXXXXXXXXXXFXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXX4 
                           => MXXXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXYXLXXXXXX1 
                           => MXXXXXXXXXXXXXXYXLXXXXXX, MXXXXXXXXXXXXXXYXLXXXX 
                           => MXXXXXXXXXXXXXXYXLXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, XFXXXXXXXXXXX => 
                           XFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXX28, 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, MXXXXXXXXXXXXXXLXXXVXX 
                           => MXXXXXXXXXXXXXXLXXXVXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1 => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, XFXXXXXXXXXXX0 => 
                           XFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, MXXXXXXXXXXXXXXXXXXMXXX
                           => MXXXXXXXXXXXXXXXXXXMXXX, 
                           MXXXXXXXXXXXXXXXXXXMXXXXX => 
                           MXXXXXXXXXXXXXXXXXXMXXXXX, MXXXXXXXXXXXXXXXXXXMXXX0 
                           => MXXXXXXXXXXXXXXXXXXMXXX1, 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, MXXXXXXXXXXXXXXXXXX0 
                           => MXXXXXXXXXXXXXXXXXX30, MXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXX31, XFXWX => sfrwe0, 
                           MXXXXXXXXXXXXXXFX => MXXXXXXXXXXXXXXFX, 
                           MXXXXXXXXXXXXXXXXXXXX6 => MXXXXXXXXXXXXXXXXXXXX22, 
                           MXXXXXXXXXXXXXXFX0 => MXXXXXXXXXXXXXXFX0, 
                           MXXXXXXXXXXXXXXXXXXXX7 => MXXXXXXXXXXXXXXXXXXXX21, 
                           MXXXXXXXXXXXXXXXXVXX => MXXXXXXXXXXXXXXXXVXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, XXMXXXXXXX => 
                           ramaddr_3, MXXXXXXXXXXXXXXXXXXMXXX1 => 
                           MXXXXXXXXXXXXXXXXXXMXXX0, XXMXXXXXXX0 => ramaddr_1, 
                           XXMXXXXXXX1 => ramaddr_0, XLXPXX => clkper, 
                           MXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXX20, XX => t0, XX0 => t1, 
                           MXXXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXXXX68, 
                           XFXXXXXX(8) => sfrdatao0_7_port, XFXXXXXX(7) => 
                           sfrdatao0_6_port, XFXXXXXX(6) => sfrdatao0_5_port, 
                           XFXXXXXX(5) => sfrdatao0_4_port, XFXXXXXX(4) => 
                           sfrdatao0_3_port, XFXXXXXX(3) => sfrdatao0_2_port, 
                           XFXXXXXX(2) => sfrdatao0_1_port, 
                           MXXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXXX69,
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXX1 => MXXXXXXXXXXXXXXXXXXXXX70,
                           MXXXXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXXXXX71,
                           MXXXXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXXXXX29)
                           ;
   XXXYXXXXXX3 : XYXX0004 port map( XLXPXX => clkper, MXXXXXXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXXXXXXX20, MXXXXXXXXXXXXXXXXXXXX
                           => MXXXXXXXXXXXXXXXXXXXX18, 
                           MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXHXFXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXXXXX0,
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXLXX, MXXXXXXXXXXXXXXLXXXVXX
                           => MXXXXXXXXXXXXXXLXXXVXX, MXXXXXXXXXXXXXXXXXXXXX =>
                           MXXXXXXXXXXXXXXXXXXXXX30, XFXXXXXXXXXX => 
                           XFXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, XFXXXXXXXXXX0 => 
                           XFXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXLXXXXXXXXXX2, MXXXXXXXXXXXXXXFXWXXX 
                           => MXXXXXXXXXXXXXXFXWXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX2, 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXXXX,
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, MXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXX4, XFXXXXXXXXXX1 => XFXXXXXXXXXX0, 
                           XXMXXXXXXX => ramaddr_6, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, XFXXXXXXXXXXX => 
                           XFXXXXXXXXXXX0, XFXXXXXXXXXXX0 => XFXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0 => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0, 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, XFXWX => sfrwe0, 
                           MXXXXXXXXXXXXXXXXVXX => MXXXXXXXXXXXXXXXXVXX, 
                           XXMXXXXXXX0 => ramaddr_3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXX28, MXXXXXXXXXXXXXXMXX => 
                           MXXXXXXXXXXXXXXMXX, MXXXXXXXXXXXXXXLXXXVX => 
                           MXXXXXXXXXXXXXXLXXXVX, MXXXXXXXXXXXXXXLXXXVX0 => 
                           MXXXXXXXXXXXXXXLXXXVX0, MXXXXXXXXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXXXXXXXXX1, XXXXX => rxd0i, 
                           MXXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXXX60,
                           XXXXX0 => rxd0o, MXXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXX61, XXXX => txd0, 
                           MXXXXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXXXXX62,
                           MXXXXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXXXXX63,
                           MXXXXXXXXXXXXXXXXXXXXX4 => MXXXXXXXXXXXXXXXXXXXXX64,
                           MXXXXXXXXXXXXXXXXXXXXX5 => MXXXXXXXXXXXXXXXXXXXXX65,
                           MXXXXXXXXXXXXXXXXXXXXX6 => MXXXXXXXXXXXXXXXXXXXXX66,
                           MXXXXXXXXXXXXXXXXXXXXX7 => MXXXXXXXXXXXXXXXXXXXXX67)
                           ;
   XXXYXXXXXX4 : XYXX0003 port map( MXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXX5, XLXXPX => clkcpu, 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXXX1, XFXXXXXXXXXX => 
                           XFXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXX21, XFXXXXXXXXXXXX => 
                           XFXXXXXXXXXXXX, MXXXXXXXXXXXXXMXMPXXXXX => 
                           MXXXXXXXXXXXXXMXMPXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, MXMXXXXXXXXXXXXX => 
                           MXMXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXX16, 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0, 
                           MXMXXXXXXXXXXXXX0 => MXMXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXPXXXXXX0, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, MXMXXXXXXXXXXXXXXXXX => 
                           MXMXXXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXXXX0 => 
                           MXMXXXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX => 
                           MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX0 => 
                           MXMXXXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXX1 => 
                           MXMXXXXXXXXXXXXX0, MXMXXXXXXXX => memdatao0_0_port, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXLXXXXXLX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX22, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, XFXXXXXXXXXX0 => 
                           XFXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, XFXXXXXXXXXX1 => 
                           XFXXXXXXXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1, XFXXXXXXXXXX2 => 
                           XFXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXX =>
                           MXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXFXXXXXXXXXXX1 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXX0 
                           => MXXXXXXXXXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXX1 
                           => MXXXXXXXXXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXX2 
                           => MXXXXXXXXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXX3 
                           => MXXXXXXXXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX10 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXX4 
                           => MXXXXXXXXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX11 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX23, MXXXXXXXXXXXXXXFXWXXX =>
                           MXXXXXXXXXXXXXXFXWXXX, MXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXMXFXXXXLXXXXXXXXXXXX, 
                           MXMXXXXXXXXXXXXXXX1 => MXMXXXXXXXXXXXXXXX18, 
                           MXMXXXXXXXXXXXXXXX2 => MXMXXXXXXXXXXXXXXX15, 
                           MXXXXXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX3, XXXXXXXXXXXX => 
                           XXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXPXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, XXXXXXX => XXXXXXX30, 
                           XFXXXXXXXXX => sfrdatao0_0_port, 
                           MXXXXXXXXXXXXXXYXXXX => MXXXXXXXXXXXXXXYXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0, MXMXXXXXXXXXXXXXXX3 
                           => MXMXXXXXXXXXXXXXXX6, XFXXXXXXXXXXX => 
                           XFXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX4 => 
                           MXMXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXXXX5 => 
                           MXMXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX0, MXMXXXXXXXXXXXXXXX6 => 
                           MXMXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX, MXMXXXXXXXXXXXXXXX7 => 
                           MXMXXXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXXXX8 => 
                           MXMXXXXXXXXXXXXXXX20, MXMXXXXXXXXXXXXXXX9 => 
                           MXMXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXMXMPXXXXXXX0 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2, MXXXXXXXXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXXXXX21, MXXXXXXXXXXXXXXXXXXXMXMPXXXX 
                           => MXXXXXXXXXXXXXXXXXXXMXMPXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXX, 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXMXMPXXXXXX, 
                           MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXYXXXXXXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXPXXXX => 
                           MXXXXXXXXXXXXXXXXXXXPXXXX, MXMXXXXXXXXXXXXXXX10 => 
                           MXMXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXXXXX14, XXMXXXXX(7) => ramdatai(7), 
                           XXMXXXXX(6) => ramdatai(6), XXMXXXXX(5) => 
                           ramdatai(5), XXMXXXXX(4) => ramdatai(4), XXMXXXXX(3)
                           => ramdatai(3), XXMXXXXX(2) => ramdatai(2), 
                           XXMXXXXX(1) => ramdatai(1), XXMXXXXX(0) => 
                           ramdatai(0), MXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXX110, MXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXX33, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2, MXXXXXXXXXXXXXXXXXX7
                           => MXXXXXXXXXXXXXXXXXX16, XXXXXXXX => XXXXXXXX25, 
                           MXXXXXXXXXXXXXXXXXX8 => MXXXXXXXXXXXXXXXXXX15, 
                           XXXXXXXX0 => XXXXXXXX24, MXXXXXXXXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXX34, MXXXXXXXXXXXXXXXXXX10 => 
                           MXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXX11 => 
                           MXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXX12 => 
                           MXXXXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXX13 => 
                           MXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXX70, MXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXX13, XXMXXXX(7) => 
                           ramaddr0_7_port, XXMXXXX(6) => ramaddr_6, XXMXXXX(5)
                           => ramaddr_5, XXMXXXX(4) => ramaddr_4, XXMXXXX(3) =>
                           ramaddr_3, XXMXXXX(2) => ramaddr_2, XXMXXXX(1) => 
                           ramaddr_1, XXMXXXX(0) => ramaddr_0, 
                           MXXXXXXXXXXXXXXYXXXX0 => MXXXXXXXXXXXXXXYXXXX2, 
                           MXXXXXXXXXXXXXXXXXXXXX1 => MXXXXXXXXXXXXXXXXXXXXX17,
                           MXXXXXXXXXXXXXXXXXVXXXXXX => 
                           MXXXXXXXXXXXXXXXXXVXXXXXX, XXXXXXXX1 => XXXXXXXX23, 
                           MXXXXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXXXXX32,
                           XXXXXXXX2 => XXXXXXXX22, MXXXXXXXXXXXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXX92, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX3, 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX10, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX5, MXXXXXXXXXXXXXXXXXXX2 
                           => MXXXXXXXXXXXXXXXXXXX45, MXXXXXXXXXXXXXXXXXXXXXXX5
                           => MXXXXXXXXXXXXXXXXXXXXXXX19, 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, 
                           MXXXXXXXXXXXXXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXXXXXX8
                           => MXXXXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXX14
                           => MXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXXXXX15 => 
                           MXXXXXXXXXXXXXXXXXX18, MXXXXXXXXXXXXXXXXXXFXWXXX => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX2, 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, MXXXXXXXXXXXXXXXXXXX3
                           => MXXXXXXXXXXXXXXXXXXX108, MXXXXXXXXXXXXXXXXXXXXX4 
                           => MXXXXXXXXXXXXXXXXXXXXX25, MXMXXXXXXXXXXXXXXX11 =>
                           MXMXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXFXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX1, 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXMWXXXXXXXXXXX, XXXXXXXXXXXXXXXX 
                           => XXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXXXXXX85, MXXXXXXXXXXXXXXXXXXFXWXXX0 
                           => MXXXXXXXXXXXXXXXXXXFXWXXX0, XFXXXXXX(8) => 
                           sfrdatao0_7_port, XFXXXXXX(7) => sfrdatao0_6_port, 
                           XFXXXXXX(6) => sfrdatao0_5_port, XFXXXXXX(5) => 
                           sfrdatao0_4_port, XFXXXXXX(4) => sfrdatao0_3_port, 
                           XFXXXXXX(3) => sfrdatao0_2_port, 
                           MXXXXXXXXXXXXXPXHXXXXXX => MXXXXXXXXXXXXXPXHXXXXXX, 
                           XXMXXXXX0(7) => ramdatao(7), XXMXXXXX0(6) => 
                           ramdatao(6), XXMXXXXX0(5) => ramdatao(5), 
                           XXMXXXXX0(4) => ramdatao(4), XXMXXXXX0(3) => 
                           ramdatao(3), XXMXXXXX0(2) => ramdatao(2), 
                           XXMXXXXX0(1) => ramdatao(1), XXMXXXXX0(0) => 
                           ramdatao(0), MXXXXXXXXXXXXXPXHXXXXXX0 => 
                           MXXXXXXXXXXXXXPXHXXXXXX0, MXXXXXXXXXXXXXPXHXXXXXX1 
                           => MXXXXXXXXXXXXXPXHXXXXXX1, 
                           MXXXXXXXXXXXXXPXHXXXXXX2 => MXXXXXXXXXXXXXPXHXXXXXX2
                           , MXXXXXXXXXXXXXPXHXXXXXX3 => 
                           MXXXXXXXXXXXXXPXHXXXXXX3, MXXXXXXXXXXXXXPXHXXXXXX4 
                           => MXXXXXXXXXXXXXPXHXXXXXX4, 
                           MXXXXXXXXXXXXXPXHXXXXXX5 => MXXXXXXXXXXXXXPXHXXXXXX6
                           , MXXXXXXXXXXXXXXXXXXX5 => MXXXXXXXXXXXXXXXXXXX49, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX11, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1 => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX5, MXXXXXXXXXXXXXPXHXXXXXX6
                           => MXXXXXXXXXXXXXPXHXXXXXX5, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX2 => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, MXXXXXXXXXXXXXXYXXXX1 =>
                           MXXXXXXXXXXXXXXYXXXX, MXXXXXXXXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXXXXXX38, XXXXXXXXXXXXXXXXXX => 
                           XXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXXXXXX100, MXXXXXXXXXXXXXXXXXXXXXX0 =>
                           MXXXXXXXXXXXXXXXXXXXXXX2, XFXXXXXXXXXXXXXXXXX => 
                           XFXXXXXXXXXXXXXXXXX, XFXXXXXXXXXXXXXXXXX0 => 
                           XFXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXX16 => 
                           MXXXXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXXX5 
                           => MXXXXXXXXXXXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXX6 => MXXXXXXXXXXXXXXXXXXXXX13,
                           MXXXXXXXXXXXXXXXMXMXMXXXX => 
                           MXXXXXXXXXXXXXXXMXMXMXXXX, MXMXXXXXXXXXXXXXXX12 => 
                           MXMXXXXXXXXXXXXXXX12, MXMXXXXXXXXXXXXXXX13 => 
                           MXMXXXXXXXXXXXXXXX7, MXMXXXXXXXXXXXXXXX14 => 
                           MXMXXXXXXXXXXXXXXX19, MXMXXXXXXXXXXXXXXX15 => 
                           MXMXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXFXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, MXXXXXXXXXXXXXXXMXXX => 
                           MXXXXXXXXXXXXXXXMXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3, 
                           MXXXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXXXX23, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10, 
                           MXXXXXXXXXXXXXXXXXX17 => MXXXXXXXXXXXXXXXXXX31, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX, 
                           MXXXXXXXXXXXXXXXMXXX0 => MXXXXXXXXXXXXXXXMXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9, 
                           MXXXXXXXXXXXXXXXXXXMXXX => MXXXXXXXXXXXXXXXXXXMXXX1,
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXPXLXXXXXX => MXXXXXXXXXXXXXPXLXXXXXX6,
                           MXXXXXXXXXXXXXPXLXXXXXX0 => MXXXXXXXXXXXXXPXLXXXXXX4
                           , MXXXXXXXXXXXXXPXLXXXXXX1 => 
                           MXXXXXXXXXXXXXPXLXXXXXX3, MXXXXXXXXXXXXXPXLXXXXXX2 
                           => MXXXXXXXXXXXXXPXLXXXXXX2, 
                           MXXXXXXXXXXXXXPXLXXXXXX3 => MXXXXXXXXXXXXXPXLXXXXXX1
                           , MXXXXXXXXXXXXXPXLXXXXXX4 => 
                           MXXXXXXXXXXXXXPXLXXXXXX0, MXXXXXXXXXXXXXPXLXXXXXX5 
                           => MXXXXXXXXXXXXXPXLXXXXXX, MXXXXXXXXXXXXXXXXXX18 =>
                           MXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXXXXXX67, MXXXXXXXXXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXXXXXX115, MXXXXXXXXXXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX14, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX13, 
                           MXXXXXXXXXXXXXXYXXXXXX => MXXXXXXXXXXXXXXYXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXX10 => MXXXXXXXXXXXXXXXXXXX72, 
                           XXMXX => ramoe, MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX1
                           => MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXXXXXXXX7 => MXXXXXXXXXXXXXXXXXXXXX21,
                           MXMXXXXXXXXXXXXXXX16 => MXMXXXXXXXXXXXXXXX, 
                           MXMXXXXXXXXXXXXXXX17 => MXMXXXXXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX6, MXXXXXXXXXXXXXXXXXXXX5
                           => MXXXXXXXXXXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX1, XFXXXXXX0(7) => 
                           sfrdatai(7), XFXXXXXX0(6) => sfrdatai(6), 
                           XFXXXXXX0(5) => sfrdatai(5), XFXXXXXX0(4) => 
                           sfrdatai(4), XFXXXXXX0(3) => sfrdatai(3), 
                           XFXXXXXX0(2) => sfrdatai(2), XFXXXXXX0(1) => 
                           sfrdatai(1), XFXXXXXX0(0) => sfrdatai(0), 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX6, XFXXXXXXXXXXX0 => 
                           XFXXXXXXXXXXX, MXXXXXXXXXXXXXXXMXXX1 => 
                           MXXXXXXXXXXXXXXXMXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX, 
                           MXXXXXXXXXXXXXXXXXX19 => MXXXXXXXXXXXXXXXXXX25, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11, 
                           MXXXXXXXXXXXXXXXXXX20 => MXXXXXXXXXXXXXXXXXX24, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX0, MXXXXXXXXXXXXXXXMXXX2 
                           => MXXXXXXXXXXXXXXXMXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXX11 => MXXXXXXXXXXXXXXXXXXX83, 
                           MXXXXXXXXXXXXXXYXXXX2 => MXXXXXXXXXXXXXXYXXXX1, 
                           MXXXXXXXXXXXXXXYXX => MXXXXXXXXXXXXXXYXX1, 
                           MXXXXXXXXXXXXXXXXXXX12 => MXXXXXXXXXXXXXXXXXXX111, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX, MXXXXXXXXXXXXXXXXXXMXXX0 
                           => MXXXXXXXXXXXXXXXXXXMXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12, 
                           MXXXXXXXXXXXXXPXLXXXXXX6 => MXXXXXXXXXXXXXPXLXXXXXX5
                           , MXXXXXXXXXXXXXXXXXX21 => MXXXXXXXXXXXXXXXXXX20, 
                           MXMXXXXXXXXXXXXXXX18 => MXMXXXXXXXXXXXXXXX0, 
                           MXMXXXXXXXXXXXXXXX19 => MXMXXXXXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXXXXX22 => MXXXXXXXXXXXXXXXXXX29, 
                           XFXWX => sfrwe0, MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4
                           => MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXX0, MXXXXXXXXXXXXXXXXXX23 
                           => MXXXXXXXXXXXXXXXXXX30, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX6, 
                           MXXXXXXXXXXXXXXXMXXX3 => MXXXXXXXXXXXXXXXMXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4, 
                           MXXXXXXXXXXXXXXXXXXMXXXXX => 
                           MXXXXXXXXXXXXXXXXXXMXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX9 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX8, 
                           MXXXXXXXXXXXXXXXXXXXHXXX => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0, MXXXXXXXXXXXXXXXXXXFXWX 
                           => MXXXXXXXXXXXXXXXXXXFXWX, MXXXXXXXXXXXXXXXMXXX4 =>
                           MXXXXXXXXXXXXXXXMXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5, 
                           MXXXXXXXXXXXXXXXXXXMXXX1 => MXXXXXXXXXXXXXXXXXXMXXX,
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXMXXVXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX10 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX11 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX7, 
                           MXXXXXXXXXXXXXXXXXXXHXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXHXXX1, MXXXXXXXXXXXXXXXMXXX5 => 
                           MXXXXXXXXXXXXXXXMXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX4, 
                           MXXXXXXXXXXXXXXXXXXXXXX1 => MXXXXXXXXXXXXXXXXXXXXXX1
                           , MXXXXXXXXXXXXXXXXXXXXXXXVXX3 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX4, MXMXXXXXXXXXXXXX2 => 
                           MXMXXXXXXXXXXXXX4, MXMXXXXXXXXXXXXX3 => 
                           MXMXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX3 
                           => MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXPXXXXXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8, 
                           MXXXXXXXXXXXXXXXXXX24 => MXXXXXXXXXXXXXXXXXX23, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXVXXXXXXX12, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXX1, MXXXXXXXXXXXXXXXMXXX6 
                           => MXXXXXXXXXXXXXXXMXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX4 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2, MXMXXXXXXXXXXXXX4 => 
                           MXMXXXXXXXXXXXXX1, MXMXXXXXXXXXXXXX5 => 
                           MXMXXXXXXXXXXXXX2, MXMXXXXXXXXXXXXX6 => 
                           MXMXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXYXX0 => 
                           MXXXXXXXXXXXXXXYXX, MXXXXXXXXXXXXXXXXXX25 => 
                           MXXXXXXXXXXXXXXXXXX28, MXXXXXXXXXXXXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXXXXXXXX9 =>
                           MXXXXXXXXXXXXXXXXXXXXX22, 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXX10 => MXXXXXXXXXXXXXXXXXXXXX3,
                           MXXXXXXXXXXXXXXXXXXXXX11 => MXXXXXXXXXXXXXXXXXXXXX24
                           , MXXXXXXXXXXXXXXXXXX26 => MXXXXXXXXXXXXXXXXXX22, 
                           MXXXXXXXXXXXXXXXXXXXXX12 => MXXXXXXXXXXXXXXXXXXXXX56
                           , MXXXXXXXXXXXXXXXXXXXXX13 => 
                           MXXXXXXXXXXXXXXXXXXXXX57, XXMWX => ramwe, XFXXX => 
                           sfroe, MXXXXXXXXXXXXXXXXXXXXX14 => 
                           MXXXXXXXXXXXXXXXXXXXXX58, MXXXXXXXXXXXXXXXXXXXXX15 
                           => MXXXXXXXXXXXXXXXXXXXXX59);
   XXXYXXXXXX5 : XYXX0002 port map( MXXXXXXXXXXXXXXXXXXXFXWXXX => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX0, MXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXX71, MXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXX14, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXXXX, XLXXPX => clkcpu, 
                           MXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXPXLXXXXXX 
                           => MXXXXXXXXXXXXXPXLXXXXXX5, ramaddr(5) => ramaddr_4
                           , ramaddr(4) => ramaddr_3, ramaddr(3) => ramaddr_2, 
                           XFXXXXXXXXXX => XFXXXXXXXXXX, XFXXXXXXXXXXXX => 
                           XFXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXFXWXXX0 => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX5, MXXXXXXXXXXXXXXYXX => 
                           MXXXXXXXXXXXXXXYXX, MXXXXXXXXXXXXXMXMPXXXXXXX => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX, MXXXXXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXXXXXX1, 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHX, 
                           MXXXXXXXXXXXXXMXMPXXXXXX => MXXXXXXXXXXXXXMXMPXXXXXX
                           , MXMPXXXXWXXX => MXMPXXXXWXXX, 
                           MXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXX66, 
                           MXXXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXXXX2
                           , MXXXXXXXXXXXXXXYXXXXXX => MXXXXXXXXXXXXXXYXXXXXX, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXXXX, MXXXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXXXX13, MXMPXXX => mempsrd, 
                           XFXXXXXXXXXX0 => XFXXXXXXXXXX0, XFXXXXXXXXXX1 => 
                           XFXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXFXWXXXXX => 
                           MXXXXXXXXXXXXXXXXXXFXWXXXXX, XXXXXPXXX => XXXXXPXXX,
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXX, MXXXXXXXXXXXXXXYXXXX 
                           => MXXXXXXXXXXXXXXYXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX, 
                           MXXXXXXXXXXXXXXXXXFXXXHX => MXXXXXXXXXXXXXXXXXFXXXHX
                           , MXXXXXXXXXXXXXXXXXXLLXX => MXXXXXXXXXXXXXXXXXXLLXX
                           , MXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXX34, MXXXXXXXXXXXXXPXLXXXXXX0 
                           => MXXXXXXXXXXXXXPXLXXXXXX4, 
                           MXXXXXXXXXXXXXPXLXXXXXX1 => MXXXXXXXXXXXXXPXLXXXXXX3
                           , MXXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXX33, MXXXXXXXXXXXXXPXLXXXXXX2 
                           => MXXXXXXXXXXXXXPXLXXXXXX2, XXXXXXXX => XXXXXXXX23,
                           MXXXXXXXXXXXXXPXLXXXXXX3 => MXXXXXXXXXXXXXPXLXXXXXX1
                           , MXXXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXX32, MXXXXXXXXXXXXXPXLXXXXXX4 
                           => MXXXXXXXXXXXXXPXLXXXXXX0, XXXXXXXX0 => XXXXXXXX22
                           , MXXXXXXXXXXXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXXXXXXXX31, MXXXXXXXXXXXXXPXHXXXXXX =>
                           MXXXXXXXXXXXXXPXHXXXXXX0, MXXXXXXXXXXXXXPXHXXXXXX0 
                           => MXXXXXXXXXXXXXPXHXXXXXX, MXMXXXX(15) => 
                           memaddr0_15_port, MXMXXXX(14) => memaddr0_14_port, 
                           MXMXXXX(13) => memaddr0_13_port, MXMXXXX(12) => 
                           memaddr0_12_port, MXMXXXX(11) => memaddr0_11_port, 
                           MXMXXXX(10) => memaddr0_10_port, MXMXXXX(9) => 
                           memaddr0_9_port, MXMXXXX(8) => memaddr0_8_port, 
                           MXMXXXX(7) => memaddr0_7_port, MXMXXXX(6) => 
                           memaddr0_6_port, MXMXXXX(5) => memaddr0_5_port, 
                           MXMXXXX(4) => memaddr0_4_port, MXMXXXX(3) => 
                           memaddr0_3_port, MXMXXXX(2) => memaddr0_2_port, 
                           MXMXXXX(1) => memaddr0_1_port, MXMXXXX(0) => 
                           memaddr0_0_port, XXXXXXXX1 => XXXXXXXX25, XXXXXXXX2 
                           => XXXXXXXX24, MXXXXXXXXXXXXXXXXVXXXXXX => 
                           MXXXXXXXXXXXXXXXXVXXXXXX3, MXXXXXXXXXXXXXXXXXXXXXXX 
                           => MXXXXXXXXXXXXXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXXXVXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXVXXXXXX2, MXXXXXXXXXXXXXXXXVXXXXXX1
                           => MXXXXXXXXXXXXXXXXVXXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX12, 
                           MXXXXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX19, 
                           MXXXXXXXXXXXXXXXXVXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXVXXXXXX3 => 
                           MXXXXXXXXXXXXXXXXVXXXXXX0, MXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXXXXXX39, MXXXXXXXXXXXXXXXXXXPXXXXXXXX
                           => MXXXXXXXXXXXXXXXXXXPXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXVXXXXXX => 
                           MXXXXXXXXXXXXXXXXXVXXXXXX, MXXXXXXXXXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXXXXXX106, MXXXXXXX => MXXXXXXX8, 
                           MXXXXXXXXXXXXXXXXXXXHXXX => 
                           MXXXXXXXXXXXXXXXXXXXHXXX0, MXXXXXXXXXXXXXXXXXXXHXXX0
                           => MXXXXXXXXXXXXXXXXXXXHXXX, 
                           MXXXXXXXXXXXXXXXXXXXHXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXHXXX1, MXXXXXXXXXXXXXXXXXXXXX4 
                           => MXXXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXX5 
                           => MXXXXXXXXXXXXXXXXXXX75, MXXXXXXXXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXXXXXX103, XXXXXXXXXXXXXXXX => 
                           XXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXXXXXX10, MXMXXXX0 => memacki, 
                           MXXXXXXXXXXXXXXXXXXX8 => MXXXXXXXXXXXXXXXXXXX45, 
                           MXXXXXXXXXXXXXXXXVXLXX => MXXXXXXXXXXXXXXXXVXLXX, 
                           MXXXXXXXXXXXXXXXXXXX9 => MXXXXXXXXXXXXXXXXXXX108, 
                           MXXXXXXXXXXXXXXXXXXX10 => MXXXXXXXXXXXXXXXXXXX95, 
                           MXXXXXXXXXXXXXXYXXXX0 => MXXXXXXXXXXXXXXYXXXX2, 
                           MXXXXXXXXXXXXXXXXXXX11 => MXXXXXXXXXXXXXXXXXXX117, 
                           MXXXXXXXXXXXXXXXXXXX12 => MXXXXXXXXXXXXXXXXXXX40, 
                           MXXXXXXXXXXXXXXXXXXX13 => MXXXXXXXXXXXXXXXXXXX41, 
                           MXXXXXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX14, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4, 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX8 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX10 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX11 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX12 => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXVXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX0, MXXXXXXXXXXXXXXFXWXXX 
                           => MXXXXXXXXXXXXXXFXWXXX, XXMXXXXX(7) => ramdatai(7)
                           , XXMXXXXX(6) => ramdatai(6), XXMXXXXX(5) => 
                           ramdatai(5), XXMXXXXX(4) => ramdatai(4), XXMXXXXX(3)
                           => ramdatai(3), XXMXXXXX(2) => ramdatai(2), 
                           XXMXXXXX(1) => ramdatai(1), XXMXXXXX(0) => 
                           ramdatai(0), MXXXXXXXXXXXXXXFXXXXXMXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXMXXXXX, MXMXXXXXXXXXXXXXXX => 
                           MXMXXXXXXXXXXXXXXX20, MXMXXXXXXXXXXXXXXX0 => 
                           MXMXXXXXXXXXXXXXXX17, MXXXXXXXXXXXXXPXHXXXXXX1 => 
                           MXXXXXXXXXXXXXPXHXXXXXX3, MXXXXXXXXXXXXXPXHXXXXXX2 
                           => MXXXXXXXXXXXXXPXHXXXXXX4, 
                           MXXXXXXXXXXXXXPXHXXXXXX3 => MXXXXXXXXXXXXXPXHXXXXXX5
                           , MXXXXXXXXXXXXXPXHXXXXXX4 => 
                           MXXXXXXXXXXXXXPXHXXXXXX6, MXXXXXXXXXXXXXPXLXXXXXX5 
                           => MXXXXXXXXXXXXXPXLXXXXXX6, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX1 => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX4, MXMXXXXXXXXXXXXXXX1 => 
                           MXMXXXXXXXXXXXXXXX11, MXMXXXXXXXXXXXXXXX2 => 
                           MXMXXXXXXXXXXXXXXX13, MXMXXXXXXXXXXXXXXX3 => 
                           MXMXXXXXXXXXXXXXXX4, MXXXXXXXXXXXXXPXHXXXXXX5 => 
                           MXXXXXXXXXXXXXPXHXXXXXX1, MXXXXXXXXXXXXXPXHXXXXXX6 
                           => MXXXXXXXXXXXXXPXHXXXXXX2, 
                           MXXXXXXXXXXXXXPXLXXXXXX6 => MXXXXXXXXXXXXXPXLXXXXXX,
                           MXXXXXXXXXXXXXXYXX0 => MXXXXXXXXXXXXXXYXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX6, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1, MXXXXXXXXXXXXXXXXXXX14 
                           => MXXXXXXXXXXXXXXXXXXX16, MXXXXXXXXXXXXXXXJXMP => 
                           MXXXXXXXXXXXXXXXJXMP, MXXXXXXXXXXXXXXXXXXX15 => 
                           MXXXXXXXXXXXXXXXXXXX101, MXXXXXXXXXXXXXXXXXMXVXWXXX 
                           => MXXXXXXXXXXXXXXXXXMXVXWXXX, 
                           MXXXXXXXXXXXXXXXXXXX16 => MXXXXXXXXXXXXXXXXXXX34, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, MXXXXXXXXXXXXXXXXXXXX0 
                           => MXXXXXXXXXXXXXXXXXXXX12, 
                           MXXXXXXXXXXXXXXXXXXFXWXXX2 => 
                           MXXXXXXXXXXXXXXXXXXFXWXXX3, 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, MXMXXXXXXXXXXXXXXX4 => 
                           MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX5 => 
                           MXMXXXXXXXXXXXXXXX6, MXMXXXXXXXXXXXXXXX6 => 
                           MXMXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXFXXXHX => 
                           MXXXXXXXXXXXXXXXXXXFXXXHX, 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX => 
                           MXXXXXXXXXXXXXXXMXMXXXLXXXXXXXXXFXXXHXXX, 
                           MXXXXXXXXXXXXXXYXXXX1 => MXXXXXXXXXXXXXXYXXXX, 
                           MXXXXXXXXXXXXXXXXXXXX1 => MXXXXXXXXXXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXXXXXX17 => MXXXXXXXXXXXXXXXXXXX83, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXXXXXLL => MXXXXXXXXXXXXXXXXXXLL, 
                           MXMXXXXX(7) => memdatao0_7_port, MXMXXXXX(6) => 
                           memdatao0_6_port, MXMXXXXX(5) => memdatao0_5_port, 
                           MXMXXXXX(4) => memdatao0_4_port, MXMXXXXX(3) => 
                           memdatao0_3_port, MXMXXXXX(2) => memdatao0_2_port, 
                           MXMXXXXX(1) => memdatao0_1_port, MXMXXXXX(0) => 
                           memdatao0_0_port, MXMXXXXXXXXXXXXXXX7 => 
                           MXMXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXXPXXXX => 
                           MXXXXXXXXXXXXXXXXXXXPXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, XFXXXXXXXXXXX => 
                           XFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXFXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXX, MXMXXXXXXXXXXXXXXX8 => 
                           MXMXXXXXXXXXXXXXXX3, MXMXXXXXXXXXXXXXXX9 => 
                           MXMXXXXXXXXXXXXXXX10, MXMXXXXXXXXXXXXXXX10 => 
                           MXMXXXXXXXXXXXXXXX16, MXMXXXXXXXXXXXXXXX11 => 
                           MXMXXXXXXXXXXXXXXX19, MXMXXXXXXXXXXXXXXX12 => 
                           MXMXXXXXXXXXXXXXXX12, MXMXXXXXXXXXXXXXXX13 => 
                           MXMXXXXXXXXXXXXXXX7, MXMXXXXXXXXXXXXXXX14 => 
                           MXMXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXX18 => 
                           MXXXXXXXXXXXXXXXXXXX102, MXXXXXXXXXXXXXXYFLXX => 
                           MXXXXXXXXXXXXXXYFLXX, MXXXXXXXXXXXXXXXXXXX19 => 
                           MXXXXXXXXXXXXXXXXXXX69, MXXXXXXXXXXXXXXYXX1 => 
                           MXXXXXXXXXXXXXXYXX1, MXXXXXXXXXXXXXXXXXXPXXLXX => 
                           MXXXXXXXXXXXXXXXXXXPXXLXX, MXXXXXXXXXXXXXXXXXXX20 =>
                           MXXXXXXXXXXXXXXXXXXX14, MXXXXXXXXXXXXXXXXXXXXXXX3 =>
                           MXXXXXXXXXXXXXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, XXXXXXXXXXXX => 
                           XXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXX9, MXMXXXXXXXXXXXXXXX15 => 
                           MXMXXXXXXXXXXXXXXX18, MXMXXXXXXXXXXXXXXX16 => 
                           MXMXXXXXXXXXXXXXXX15, MXMXXXXXXXXXXXXX => 
                           MXMXXXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX0, XFXWX => sfrwe0, 
                           MXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXX20, 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX => 
                           MXXXXXXXXXXXXXXXXXXMXMPXXXX, MXXXXXXXXXXXXXXXXXXX21 
                           => MXXXXXXXXXXXXXXXXXXX107, XXMXXXXXXX => ramaddr_0,
                           MXXXXXXXXXXXXXMXMPXXXXX => MXXXXXXXXXXXXXMXMPXXXXX, 
                           XXXXXXXX3 => XXXXXXXX26, MXXXXXXXXXXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXXXXXXX24, MXXXXXXXXXXXXXXXXXFXXXHXXX 
                           => MXXXXXXXXXXXXXXXXXFXXXHXXX, MXXXXXXXXXXXXXXXXXX0 
                           => MXXXXXXXXXXXXXXXXXX22, MXMXXXXXXXXXXXXX0 => 
                           MXMXXXXXXXXXXXXX3, MXXXXXXXXXXXXXXFXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXX1 =>
                           MXXXXXXXXXXXXXXXXXX28, MXXXXXXXXXXXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXXXXXXXX41, MXXXXXXXXXXXXXXXXXXXXX6 =>
                           MXXXXXXXXXXXXXXXXXXXXX53, MXXXXXXXXXXXXXXXMXMXMXXXX 
                           => MXXXXXXXXXXXXXXXMXMXMXXXX, 
                           MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF => 
                           MXXXXXXXXXXXXXXXMXMXXXLXFLXXHXFF, MXMWXXXXXX => 
                           MXMWXXXXXX0, MXXXXXXXXXXXXXMXMXXXX => 
                           MXXXXXXXXXXXXXMXMXXXX, MXMXX => memrd, XFXXXXXX(7) 
                           => sfrdatao0_7_port, XFXXXXXX(6) => sfrdatao0_6_port
                           , XFXXXXXX(5) => sfrdatao0_5_port, XFXXXXXX(4) => 
                           sfrdatao0_4_port, XFXXXXXX(3) => sfrdatao0_3_port, 
                           XFXXXXXX(2) => sfrdatao0_2_port, XFXXXXXX(1) => 
                           sfrdatao0_1_port, XFXXXXXX(0) => sfrdatao0_0_port, 
                           MXXXXXXXXXXXXXXXXXXXXX7 => MXXXXXXXXXXXXXXXXXXXXX52,
                           MXMXXXXXXXXXXXXX1 => MXMXXXXXXXXXXXXX0, 
                           MXMXXXXXXXXXXXXX2 => MXMXXXXXXXXXXXXX6, 
                           MXMXXXXXXXXXXXXX3 => MXMXXXXXXXXXXXXX5, 
                           MXMXXXXXXXXXXXXX4 => MXMXXXXXXXXXXXXX4, 
                           MXMXXXXXXXXXXXXX5 => MXMXXXXXXXXXXXXX1, 
                           MXMXXXXXXXXXXXXX6 => MXMXXXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXXXX8 => MXXXXXXXXXXXXXXXXXXXXX51,
                           MXXXXXXXXXXXXXXXXXXXXX9 => MXXXXXXXXXXXXXXXXXXXXX50,
                           MXXXXXXXXXXXXXXXXXXXXX10 => MXXXXXXXXXXXXXXXXXXXXX49
                           , MXXXXXXXXXXXXXXXXXXXXX11 => 
                           MXXXXXXXXXXXXXXXXXXXXX48, MXXXXXXXXXXXXXXXXXXXXX12 
                           => MXXXXXXXXXXXXXXXXXXXXX47, 
                           MXXXXXXXXXXXXXXXXXXXXX13 => MXXXXXXXXXXXXXXXXXXXXX46
                           , MXXXXXXXXXXXXXXXXXXXXX14 => 
                           MXXXXXXXXXXXXXXXXXXXXX45);
   XXXYXXXXXX6 : XYXX0001 port map( MXXXXXXXXXXXXXMXMXXXX => 
                           MXXXXXXXXXXXXXMXMXXXX, XLXXPX => clkcpu, 
                           MXXXXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXXXXX4,
                           MXXXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXXXX34, 
                           XXXXXXXX => XXXXXXXX25, MXXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXX3, XXXXXXXX0 => XXXXXXXX24, 
                           MXXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXXX33,
                           XXXXXXXX1 => XXXXXXXX23, MXXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXX32, XXXXXXXX2 => XXXXXXXX22, 
                           MXXXXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXXXXX31,
                           MXXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXXX15, 
                           MXMXXXXXXXXXXXXX => MXMXXXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXX17, 
                           MXXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXXX14, 
                           MXXXXXXXXXXXXXXXXXXX => MXXXXXXXXXXXXXXXXXXX57, 
                           MXXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXXX8, 
                           MXXXXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXXXXX27,
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXX15, 
                           MXXXXXXXXXXXXXXXXXX0 => MXXXXXXXXXXXXXXXXXX16, 
                           MXXXXXXXXXXXXXXXXXX1 => MXXXXXXXXXXXXXXXXXX15, 
                           MXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXX14, 
                           MXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXX13, 
                           MXXXXXXXXXXXXXXXXXX4 => MXXXXXXXXXXXXXXXXXX12, 
                           MXXXXXXXXXXXXXXFXWXXX => MXXXXXXXXXXXXXXFXWXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX1, MXXXXXXXXXXXXXXYXX => 
                           MXXXXXXXXXXXXXXYXX0, MXXXXXXXXXXXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXX15, MXXXXXXXXXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXX123, MXXXXXXXXXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXFXWXXXXX 
                           => MXXXXXXXXXXXXXXXXXXFXWXXXXX, XFXXXXXXXXXX => 
                           XFXXXXXXXXXX2, XFXXXXXXXXXX0 => XFXXXXXXXXXX, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX1, MXXXXXXXXXXXXXXXXXXX4 
                           => MXXXXXXXXXXXXXXXXXXX93, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX1, MXXXXXXXXXXXXXXXXXXX5 
                           => MXXXXXXXXXXXXXXXXXXX118, MXXXXXXXXXXXXXXXXXXX6 =>
                           MXXXXXXXXXXXXXXXXXXX71, MXXXXXXXXXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXXXXXX66, MXXXXXXXXXXXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXXXXXX119, XFXXXXXXXXXXX => 
                           XFXXXXXXXXXXX0, MXXXXXXXXXXXXXXFXXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXX4, MXXXXXXXXXXXXXXXXXXX9 
                           => MXXXXXXXXXXXXXXXXXXX65, MXXXXXXXXXXXXXXXXXXX10 =>
                           MXXXXXXXXXXXXXXXXXXX116, MXXXXXXXXXXXXXXXXXXX11 => 
                           MXXXXXXXXXXXXXXXXXXX109, MXXXXXXXXXXXXXXXXXXX12 => 
                           MXXXXXXXXXXXXXXXXXXX63, MXXXXXXXXXXXXXXXXXXX13 => 
                           MXXXXXXXXXXXXXXXXXXX87, MXXXXXXXXXXXXXMXMPXXXXXXX0 
                           => MXXXXXXXXXXXXXMXMPXXXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXX14 => MXXXXXXXXXXXXXXXXXXX89, 
                           MXXXXXXXXXXXXXXXXXXXXX6 => MXXXXXXXXXXXXXXXXXXXXX20,
                           MXXXXXXXXXXXXXXXXXXX15 => MXXXXXXXXXXXXXXXXXXX86, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXX16 => MXXXXXXXXXXXXXXXXXXX61, 
                           MXXXXXXXXXXXXXXXXXXX17 => MXXXXXXXXXXXXXXXXXXX104, 
                           MXXXXXXXXXXXXXXXXXXX18 => MXXXXXXXXXXXXXXXXXXX84, 
                           MXXXXXXXXXXXXXXXXXXX19 => MXXXXXXXXXXXXXXXXXXX91, 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXVXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXX7 => MXXXXXXXXXXXXXXXXXXXXX15,
                           MXXXXXXXXXXXXXXXXXXXXX8 => MXXXXXXXXXXXXXXXXXXXXX14,
                           MXXXXXXXXXXXXXXXXXXX20 => MXXXXXXXXXXXXXXXXXXX14, 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX, MXXXXXXXXXXXXXXYXXXX => 
                           MXXXXXXXXXXXXXXYXXXX2, MXXXXXXXXXXXXXXXXXXX21 => 
                           MXXXXXXXXXXXXXXXXXXX38, 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX => 
                           MXXXXXXXXXXXXXXXXXPXWXXXXWXXX, XFXXXXXXXXXX1 => 
                           XFXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXFXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXFXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXX1, MXXXXXXXXXXXXXXYXXXX0 => 
                           MXXXXXXXXXXXXXXYXXXX1, MXXXXXXXXXXXXXXFXXXXXXXXXX =>
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX1 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX5 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX3, 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX6 => 
                           MXXXXXXXXXXXXXXFXXXXXXLXXXVXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXX22 => MXXXXXXXXXXXXXXXXXXX7, 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX => 
                           MXXXXXXXXXXXXXXXXXXXFXWXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX3, MXXXXXXXXXXXXXXXXXXX23
                           => MXXXXXXXXXXXXXXXXXXX88, 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXPXXXXXXXX, MXXXXXXXXXXXXXXYXXXX1 
                           => MXXXXXXXXXXXXXXYXXXX0, MXXXXXXXXXXXXXXXXXXX24 => 
                           MXXXXXXXXXXXXXXXXXXX0, MXXXXXXXXXXXXXXXXXXX25 => 
                           MXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXX26 => 
                           MXXXXXXXXXXXXXXXXXXX120, MXXXXXXXXXXXXXXXXXXX27 => 
                           MXXXXXXXXXXXXXXXXXXX50, MXXXXXXXXXXXXXXXXXXX28 => 
                           MXXXXXXXXXXXXXXXXXXX90, MXXXXXXXXXXXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXX29 => 
                           MXXXXXXXXXXXXXXXXXXX82, MXXXXXXXXXXXXXXXXXX5 => 
                           MXXXXXXXXXXXXXXXXXX11, MXXXXXXXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXXXXX10, MXXXXXXXXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXX8 => 
                           MXXXXXXXXXXXXXXXXXX8, MXXXXXXXXXXXXXXXXXX9 => 
                           MXXXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXXXXX10 => 
                           MXXXXXXXXXXXXXXXXXX6, MXXXXXXXXXXXXXXXXXXX30 => 
                           MXXXXXXXXXXXXXXXXXXX22, MXXXXXXXXXXXXXXXXXXXXXXXVXX0
                           => MXXXXXXXXXXXXXXXXXXXXXXXVXX8, 
                           MXXXXXXXXXXXXXXXXXX11 => MXXXXXXXXXXXXXXXXXX5, 
                           MXMXXXXXXXXXXXXXXX => MXMXXXXXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXXXXX12 => MXXXXXXXXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXXXXX13 => MXXXXXXXXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXXXXX14 => MXXXXXXXXXXXXXXXXXX2, 
                           MXMXXXXXXXXXXXXXXX0 => MXMXXXXXXXXXXXXXXX20, 
                           MXMXXXXXXXXXXXXXXX1 => MXMXXXXXXXXXXXXXXX16, 
                           MXMXXXXXXXXXXXXXXX2 => MXMXXXXXXXXXXXXXXX1, 
                           MXMXXXXXXXXXXXXXXX3 => MXMXXXXXXXXXXXXXXX9, 
                           MXMXXXXXXXXXXXXXXX4 => MXMXXXXXXXXXXXXXXX11, 
                           MXMXXXXXXXXXXXXXXX5 => MXMXXXXXXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXXXXXX31 => MXXXXXXXXXXXXXXXXXXX80, 
                           MXXXXXXXXXXXXXXYXXXX2 => MXXXXXXXXXXXXXXYXXXX, 
                           MXXXXXXXXXXXXXMXMPXXXXXXX1 => 
                           MXXXXXXXXXXXXXMXMPXXXXXXX0, MXXXXXXXXXXXXXXXXXXXX2 
                           => MXXXXXXXXXXXXXXXXXXXX12, MXXXXXXXXXXXXXXXXXXX32 
                           => MXXXXXXXXXXXXXXXXXXX34, MXXXXXXX => MXXXXXXX4, 
                           MXXXXXXXXXXXXXXXXLXXXXXXX => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX0, 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX => 
                           MXXXXXXXXXXXXXXXXLXXXLXXXXXLXXXVXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXX10 => MXXXXXXXXXXXXXXXXXXXXX12
                           , MXXXXXXXXXXXXXXXXXXXXX11 => 
                           MXXXXXXXXXXXXXXXXXXXXX9, MXXXXXXXXXXXXXXXXXXXXXX1 =>
                           MXXXXXXXXXXXXXXXXXXXXXX2, MXXXXXXXXXXXXXXXXXXXXXVXX 
                           => MXXXXXXXXXXXXXXXXXXXXXVXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXX0, MXXXXXXXXXXXXXXXXXXX33 
                           => MXXXXXXXXXXXXXXXXXXX122, 
                           MXXXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXX15, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXYFLXX => 
                           MXXXXXXXXXXXXXXYFLXX, MXXXXXXXXXXXXXXXXXXXXX12 => 
                           MXXXXXXXXXXXXXXXXXXXXX8, MXMXXXXX(7) => 
                           memdatao0_7_port, MXMXXXXX(6) => memdatao0_6_port, 
                           MXMXXXXX(5) => memdatao0_5_port, MXMXXXXX(4) => 
                           memdatao0_4_port, MXMXXXXX(3) => memdatao0_3_port, 
                           MXMXXXXX(2) => memdatao0_2_port, MXMXXXXX(1) => 
                           memdatao0_1_port, MXMXXXXX(0) => memdatao0_0_port, 
                           MXXXXXXXXXXXXXXXXXXXX3 => MXXXXXXXXXXXXXXXXXXXX11, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX5, 
                           MXXXXXXXXXXXXXXXXXXXXX13 => MXXXXXXXXXXXXXXXXXXXXX7,
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4, MXXXXXXXXXXXXXXXMXXX =>
                           MXXXXXXXXXXXXXXXMXXX6, MXXXXXXXXXXXXXXFXXXXXXXXXX1 
                           => MXXXXXXXXXXXXXXFXXXXXXXXXX1, 
                           MXXXXXXXXXXXXXXXMXXX0 => MXXXXXXXXXXXXXXXMXXX5, 
                           MXXXXXXXXXXXXXXXMXXX1 => MXXXXXXXXXXXXXXXMXXX4, 
                           MXXXXXXXXXXXXXXXMXXX2 => MXXXXXXXXXXXXXXXMXXX3, 
                           MXMXXXXXXXXXXXXXXX6 => MXMXXXXXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX6, MXMXXXXXXXXXXXXXXX7 
                           => MXMXXXXXXXXXXXXXXX10, MXMXXXXXXXXXXXXXXX8 => 
                           MXMXXXXXXXXXXXXXXX5, MXMXXXXXXXXXXXXXXX9 => 
                           MXMXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXXXX10 => 
                           MXMXXXXXXXXXXXXXXX19, MXXXXXXXXXXXXXXXXXXX34 => 
                           MXXXXXXXXXXXXXXXXXXX5, MXXXXXXXXXXXXXXXXXXX35 => 
                           MXXXXXXXXXXXXXXXXXXX48, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXX14 => MXXXXXXXXXXXXXXXXXXXXX6,
                           MXXXXXXXXXXXXXXXXXXXX4 => MXXXXXXXXXXXXXXXXXXXX10, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXX1, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX0, 
                           MXXXXXXXXXXXXXXXXXXXXX15 => MXXXXXXXXXXXXXXXXXXXXX0,
                           MXXXXXXXXXXXXXXXXLXXXXXXX0 => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX2, MXXXXXXXXXXXXXXXXXXX36 
                           => MXXXXXXXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXX37 => 
                           MXXXXXXXXXXXXXXXXXXX77, MXMXXXXXXXXXXXXXXX11 => 
                           MXMXXXXXXXXXXXXXXX13, MXXXXXXXXXXXXXXXXXXXXX16 => 
                           MXXXXXXXXXXXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX2 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX7, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXXXXXX1, 
                           MXXXXXXXXXXXXXXXXXXX38 => MXXXXXXXXXXXXXXXXXXX39, 
                           MXXXXXXXXXXXXXXXXXXX39 => MXXXXXXXXXXXXXXXXXXX68, 
                           MXXXXXXXXXXXXXXXXXXX40 => MXXXXXXXXXXXXXXXXXXX74, 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX3 => 
                           MXXXXXXXXXXXXXXXXXXXXXXXVXX9, MXXXXXXXXXXXXXXXXXXXX5
                           => MXXXXXXXXXXXXXXXXXXXX9, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX2 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX3, MXXXXXXXXXXXXXXXMXXX3 
                           => MXXXXXXXXXXXXXXXMXXX2, XFXXXXXXXXXXX0 => 
                           XFXXXXXXXXXXX, MXXXXXXXXXXXXXXFXXXXXXXXXX3 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX0, 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX4 => 
                           MXXXXXXXXXXXXXXFXXXXXXXXXX, ramaddr(6) => ramaddr_5,
                           ramaddr(5) => ramaddr_4, ramaddr(4) => ramaddr_3, 
                           ramaddr(3) => ramaddr_2, ramaddr(2) => ramaddr_1, 
                           ramaddr(1) => ramaddr_0, MXXXXXXXXXXXXXXXMXXX4 => 
                           MXXXXXXXXXXXXXXXMXXX0, MXXXXXXXXXXXXXXXMXXX5 => 
                           MXXXXXXXXXXXXXXXMXXX, MXXXXXXXXXXXXXXYXXXXXX => 
                           MXXXXXXXXXXXXXXYXXXXXX, MXXXXXXXXXXXXXMXMPXXXXXXX2 
                           => MXXXXXXXXXXXXXMXMPXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXX2 => MXXXXXXXXXXXXXXXXXXXXXX1
                           , MXXXXXXXXXXXXXXYXX0 => MXXXXXXXXXXXXXXYXX, 
                           MXXXXXXXXXXXXXXXXXVXXXXXX => 
                           MXXXXXXXXXXXXXXXXXVXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX0 => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX0, 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX1 => 
                           MXXXXXXXXXXXXXXXXXXXXXXWXXX, MXXXXXXXXXXXXXXXMXXX6 
                           => MXXXXXXXXXXXXXXXMXXX1, MXXXXXXXXXXXXXXXJXMP => 
                           MXXXXXXXXXXXXXXXJXMP, MXXXXXXXXXXXXXXXXVXLXX => 
                           MXXXXXXXXXXXXXXXXVXLXX, MXXXXXXXXXXXXXXXXXXXX6 => 
                           MXXXXXXXXXXXXXXXXXXXX8, MXMXXXXXXXXXXXXX0 => 
                           MXMXXXXXXXXXXXXX6, MXMXXXXXXXXXXXXX1 => 
                           MXMXXXXXXXXXXXXX, MXXXXXXXXXXXXXXXXXXXX7 => 
                           MXXXXXXXXXXXXXXXXXXXX7, MXXXXXXXXXXXXXXFXXXXXXXXXXX6
                           => MXXXXXXXXXXXXXXFXXXXXXXXXXX, 
                           MXXXXXXXXXXXXXXXXXXXX8 => MXXXXXXXXXXXXXXXXXXXX6, 
                           MXXXXXXXXXXXXXXXXXXXX9 => MXXXXXXXXXXXXXXXXXXXX5, 
                           MXXXXXXXXXXXXXXXXXXXX10 => MXXXXXXXXXXXXXXXXXXXX4, 
                           MXXXXXXXXXXXXXXXXLXXXXXXX1 => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX1, MXXXXXXXXXXXXXXXXXXXX11 
                           => MXXXXXXXXXXXXXXXXXXXX3, 
                           MXXXXXXXXXXXXXXXXLXXXXXXX2 => 
                           MXXXXXXXXXXXXXXXXLXXXXXXX, MXXXXXXXXXXXXXXXXXXXX12 
                           => MXXXXXXXXXXXXXXXXXXXX2, 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX => 
                           MXXXXXXXXXXXXXXXXXXXXXXVXXXXXXXXXXXXXXXXXXXXXXXX4);

end SYN_verilog;
